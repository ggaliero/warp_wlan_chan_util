--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_2fe7f24afe1bc972.vhd when simulating
-- the core, addsb_11_0_2fe7f24afe1bc972. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_2fe7f24afe1bc972 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END addsb_11_0_2fe7f24afe1bc972;

ARCHITECTURE addsb_11_0_2fe7f24afe1bc972_a OF addsb_11_0_2fe7f24afe1bc972 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_2fe7f24afe1bc972
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_2fe7f24afe1bc972 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 5,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "00000",
      c_b_width => 5,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 5,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_2fe7f24afe1bc972
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_2fe7f24afe1bc972_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_5c670787eb4ba225.vhd when simulating
-- the core, addsb_11_0_5c670787eb4ba225. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_5c670787eb4ba225 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END addsb_11_0_5c670787eb4ba225;

ARCHITECTURE addsb_11_0_5c670787eb4ba225_a OF addsb_11_0_5c670787eb4ba225 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_5c670787eb4ba225
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_5c670787eb4ba225 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 3,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "000",
      c_b_width => 3,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 3,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_5c670787eb4ba225
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_5c670787eb4ba225_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_60fd3b5996582b7a.vhd when simulating
-- the core, addsb_11_0_60fd3b5996582b7a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_60fd3b5996582b7a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END addsb_11_0_60fd3b5996582b7a;

ARCHITECTURE addsb_11_0_60fd3b5996582b7a_a OF addsb_11_0_60fd3b5996582b7a IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_60fd3b5996582b7a
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_60fd3b5996582b7a USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 9,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "000000000",
      c_b_width => 9,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 9,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_60fd3b5996582b7a
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_60fd3b5996582b7a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_6695c8a33176d3c2.vhd when simulating
-- the core, addsb_11_0_6695c8a33176d3c2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_6695c8a33176d3c2 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END addsb_11_0_6695c8a33176d3c2;

ARCHITECTURE addsb_11_0_6695c8a33176d3c2_a OF addsb_11_0_6695c8a33176d3c2 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_6695c8a33176d3c2
  PORT (
    a : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_6695c8a33176d3c2 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 18,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000",
      c_b_width => 18,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 18,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_6695c8a33176d3c2
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_6695c8a33176d3c2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_73986f767e994888.vhd when simulating
-- the core, addsb_11_0_73986f767e994888. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_73986f767e994888 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END addsb_11_0_73986f767e994888;

ARCHITECTURE addsb_11_0_73986f767e994888_a OF addsb_11_0_73986f767e994888 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_73986f767e994888
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_73986f767e994888 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 10,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "0000000000",
      c_b_width => 10,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 10,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_73986f767e994888
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_73986f767e994888_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_7925f33378f00f6a.vhd when simulating
-- the core, addsb_11_0_7925f33378f00f6a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_7925f33378f00f6a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END addsb_11_0_7925f33378f00f6a;

ARCHITECTURE addsb_11_0_7925f33378f00f6a_a OF addsb_11_0_7925f33378f00f6a IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_7925f33378f00f6a
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_7925f33378f00f6a USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 3,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000",
      c_b_width => 3,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 3,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_7925f33378f00f6a
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_7925f33378f00f6a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_7cf14debcedb76ce.vhd when simulating
-- the core, addsb_11_0_7cf14debcedb76ce. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_7cf14debcedb76ce IS
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END addsb_11_0_7cf14debcedb76ce;

ARCHITECTURE addsb_11_0_7cf14debcedb76ce_a OF addsb_11_0_7cf14debcedb76ce IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_7cf14debcedb76ce
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_7cf14debcedb76ce USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 13,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "0000000000000",
      c_b_width => 13,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 13,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_7cf14debcedb76ce
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_7cf14debcedb76ce_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_8942e2ad5d8d4897.vhd when simulating
-- the core, addsb_11_0_8942e2ad5d8d4897. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_8942e2ad5d8d4897 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END addsb_11_0_8942e2ad5d8d4897;

ARCHITECTURE addsb_11_0_8942e2ad5d8d4897_a OF addsb_11_0_8942e2ad5d8d4897 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_8942e2ad5d8d4897
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_8942e2ad5d8d4897 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 9,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000",
      c_b_width => 9,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 9,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_8942e2ad5d8d4897
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_8942e2ad5d8d4897_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_a52ead9b8a3c1e76.vhd when simulating
-- the core, addsb_11_0_a52ead9b8a3c1e76. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_a52ead9b8a3c1e76 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END addsb_11_0_a52ead9b8a3c1e76;

ARCHITECTURE addsb_11_0_a52ead9b8a3c1e76_a OF addsb_11_0_a52ead9b8a3c1e76 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_a52ead9b8a3c1e76
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_a52ead9b8a3c1e76 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 9,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000",
      c_b_width => 9,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 9,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_a52ead9b8a3c1e76
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_a52ead9b8a3c1e76_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_d5bf78f2384e976c.vhd when simulating
-- the core, addsb_11_0_d5bf78f2384e976c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_d5bf78f2384e976c IS
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END addsb_11_0_d5bf78f2384e976c;

ARCHITECTURE addsb_11_0_d5bf78f2384e976c_a OF addsb_11_0_d5bf78f2384e976c IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_d5bf78f2384e976c
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_d5bf78f2384e976c USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 10,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000",
      c_b_width => 10,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 10,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_d5bf78f2384e976c
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_d5bf78f2384e976c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_f66fe30ee2d0a6f0.vhd when simulating
-- the core, addsb_11_0_f66fe30ee2d0a6f0. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_f66fe30ee2d0a6f0 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(16 DOWNTO 0)
  );
END addsb_11_0_f66fe30ee2d0a6f0;

ARCHITECTURE addsb_11_0_f66fe30ee2d0a6f0_a OF addsb_11_0_f66fe30ee2d0a6f0 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_f66fe30ee2d0a6f0
  PORT (
    a : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(16 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_f66fe30ee2d0a6f0 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 17,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "00000000000000000",
      c_b_width => 17,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 17,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_f66fe30ee2d0a6f0
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_f66fe30ee2d0a6f0_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file axififo_fg92_83e0abc99b742965.vhd when simulating
-- the core, axififo_fg92_83e0abc99b742965. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY axififo_fg92_83e0abc99b742965 IS
  PORT (
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    s_axis_tuser : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    m_axis_tuser : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    axis_data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END axififo_fg92_83e0abc99b742965;

ARCHITECTURE axififo_fg92_83e0abc99b742965_a OF axififo_fg92_83e0abc99b742965 IS
-- synthesis translate_off
COMPONENT wrapped_axififo_fg92_83e0abc99b742965
  PORT (
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    s_axis_tuser : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    m_axis_tuser : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    axis_data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_axififo_fg92_83e0abc99b742965 USE ENTITY XilinxCoreLib.fifo_generator_v9_3(behavioral)
    GENERIC MAP (
      c_add_ngc_constraint => 0,
      c_application_type_axis => 0,
      c_application_type_rach => 0,
      c_application_type_rdch => 0,
      c_application_type_wach => 0,
      c_application_type_wdch => 0,
      c_application_type_wrch => 0,
      c_axi_addr_width => 32,
      c_axi_aruser_width => 1,
      c_axi_awuser_width => 1,
      c_axi_buser_width => 1,
      c_axi_data_width => 64,
      c_axi_id_width => 4,
      c_axi_ruser_width => 1,
      c_axi_type => 0,
      c_axi_wuser_width => 1,
      c_axis_tdata_width => 32,
      c_axis_tdest_width => 4,
      c_axis_tid_width => 8,
      c_axis_tkeep_width => 4,
      c_axis_tstrb_width => 4,
      c_axis_tuser_width => 18,
      c_axis_type => 0,
      c_common_clock => 1,
      c_count_type => 0,
      c_data_count_width => 10,
      c_default_value => "BlankString",
      c_din_width => 18,
      c_din_width_axis => 51,
      c_din_width_rach => 32,
      c_din_width_rdch => 64,
      c_din_width_wach => 32,
      c_din_width_wdch => 64,
      c_din_width_wrch => 2,
      c_dout_rst_val => "0",
      c_dout_width => 18,
      c_enable_rlocs => 0,
      c_enable_rst_sync => 1,
      c_error_injection_type => 0,
      c_error_injection_type_axis => 0,
      c_error_injection_type_rach => 0,
      c_error_injection_type_rdch => 0,
      c_error_injection_type_wach => 0,
      c_error_injection_type_wdch => 0,
      c_error_injection_type_wrch => 0,
      c_family => "virtex6",
      c_full_flags_rst_val => 1,
      c_has_almost_empty => 0,
      c_has_almost_full => 0,
      c_has_axi_aruser => 0,
      c_has_axi_awuser => 0,
      c_has_axi_buser => 0,
      c_has_axi_rd_channel => 0,
      c_has_axi_ruser => 0,
      c_has_axi_wr_channel => 0,
      c_has_axi_wuser => 0,
      c_has_axis_tdata => 1,
      c_has_axis_tdest => 0,
      c_has_axis_tid => 0,
      c_has_axis_tkeep => 0,
      c_has_axis_tlast => 1,
      c_has_axis_tready => 1,
      c_has_axis_tstrb => 0,
      c_has_axis_tuser => 1,
      c_has_backup => 0,
      c_has_data_count => 0,
      c_has_data_counts_axis => 1,
      c_has_data_counts_rach => 0,
      c_has_data_counts_rdch => 0,
      c_has_data_counts_wach => 0,
      c_has_data_counts_wdch => 0,
      c_has_data_counts_wrch => 0,
      c_has_int_clk => 0,
      c_has_master_ce => 0,
      c_has_meminit_file => 0,
      c_has_overflow => 0,
      c_has_prog_flags_axis => 0,
      c_has_prog_flags_rach => 0,
      c_has_prog_flags_rdch => 0,
      c_has_prog_flags_wach => 0,
      c_has_prog_flags_wdch => 0,
      c_has_prog_flags_wrch => 0,
      c_has_rd_data_count => 0,
      c_has_rd_rst => 0,
      c_has_rst => 1,
      c_has_slave_ce => 0,
      c_has_srst => 0,
      c_has_underflow => 0,
      c_has_valid => 0,
      c_has_wr_ack => 0,
      c_has_wr_data_count => 0,
      c_has_wr_rst => 0,
      c_implementation_type => 0,
      c_implementation_type_axis => 1,
      c_implementation_type_rach => 2,
      c_implementation_type_rdch => 1,
      c_implementation_type_wach => 2,
      c_implementation_type_wdch => 1,
      c_implementation_type_wrch => 2,
      c_init_wr_pntr_val => 0,
      c_interface_type => 1,
      c_memory_type => 1,
      c_mif_file_name => "BlankString",
      c_msgon_val => 1,
      c_optimization_mode => 0,
      c_overflow_low => 0,
      c_preload_latency => 1,
      c_preload_regs => 0,
      c_prim_fifo_type => "4kx4",
      c_prog_empty_thresh_assert_val => 2,
      c_prog_empty_thresh_assert_val_axis => 126,
      c_prog_empty_thresh_assert_val_rach => 14,
      c_prog_empty_thresh_assert_val_rdch => 1022,
      c_prog_empty_thresh_assert_val_wach => 14,
      c_prog_empty_thresh_assert_val_wdch => 1022,
      c_prog_empty_thresh_assert_val_wrch => 14,
      c_prog_empty_thresh_negate_val => 3,
      c_prog_empty_type => 0,
      c_prog_empty_type_axis => 0,
      c_prog_empty_type_rach => 0,
      c_prog_empty_type_rdch => 0,
      c_prog_empty_type_wach => 0,
      c_prog_empty_type_wdch => 0,
      c_prog_empty_type_wrch => 0,
      c_prog_full_thresh_assert_val => 1022,
      c_prog_full_thresh_assert_val_axis => 127,
      c_prog_full_thresh_assert_val_rach => 15,
      c_prog_full_thresh_assert_val_rdch => 1023,
      c_prog_full_thresh_assert_val_wach => 15,
      c_prog_full_thresh_assert_val_wdch => 1023,
      c_prog_full_thresh_assert_val_wrch => 15,
      c_prog_full_thresh_negate_val => 1021,
      c_prog_full_type => 0,
      c_prog_full_type_axis => 0,
      c_prog_full_type_rach => 0,
      c_prog_full_type_rdch => 0,
      c_prog_full_type_wach => 0,
      c_prog_full_type_wdch => 0,
      c_prog_full_type_wrch => 0,
      c_rach_type => 0,
      c_rd_data_count_width => 10,
      c_rd_depth => 1024,
      c_rd_freq => 1,
      c_rd_pntr_width => 10,
      c_rdch_type => 0,
      c_reg_slice_mode_axis => 0,
      c_reg_slice_mode_rach => 0,
      c_reg_slice_mode_rdch => 0,
      c_reg_slice_mode_wach => 0,
      c_reg_slice_mode_wdch => 0,
      c_reg_slice_mode_wrch => 0,
      c_synchronizer_stage => 2,
      c_underflow_low => 0,
      c_use_common_overflow => 0,
      c_use_common_underflow => 0,
      c_use_default_settings => 0,
      c_use_dout_rst => 1,
      c_use_ecc => 0,
      c_use_ecc_axis => 0,
      c_use_ecc_rach => 0,
      c_use_ecc_rdch => 0,
      c_use_ecc_wach => 0,
      c_use_ecc_wdch => 0,
      c_use_ecc_wrch => 0,
      c_use_embedded_reg => 0,
      c_use_fifo16_flags => 0,
      c_use_fwft_data_count => 0,
      c_valid_low => 0,
      c_wach_type => 0,
      c_wdch_type => 0,
      c_wr_ack_low => 0,
      c_wr_data_count_width => 10,
      c_wr_depth => 1024,
      c_wr_depth_axis => 128,
      c_wr_depth_rach => 16,
      c_wr_depth_rdch => 1024,
      c_wr_depth_wach => 16,
      c_wr_depth_wdch => 1024,
      c_wr_depth_wrch => 16,
      c_wr_freq => 1,
      c_wr_pntr_width => 10,
      c_wr_pntr_width_axis => 7,
      c_wr_pntr_width_rach => 4,
      c_wr_pntr_width_rdch => 10,
      c_wr_pntr_width_wach => 4,
      c_wr_pntr_width_wdch => 10,
      c_wr_pntr_width_wrch => 4,
      c_wr_response_latency => 1,
      c_wrch_type => 0
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_axififo_fg92_83e0abc99b742965
  PORT MAP (
    s_aclk => s_aclk,
    s_aresetn => s_aresetn,
    s_axis_tvalid => s_axis_tvalid,
    s_axis_tready => s_axis_tready,
    s_axis_tdata => s_axis_tdata,
    s_axis_tlast => s_axis_tlast,
    s_axis_tuser => s_axis_tuser,
    m_axis_tvalid => m_axis_tvalid,
    m_axis_tready => m_axis_tready,
    m_axis_tdata => m_axis_tdata,
    m_axis_tlast => m_axis_tlast,
    m_axis_tuser => m_axis_tuser,
    axis_data_count => axis_data_count
  );
-- synthesis translate_on

END axififo_fg92_83e0abc99b742965_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_30fab105208816ae.vhd when simulating
-- the core, bmg_72_30fab105208816ae. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_30fab105208816ae IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END bmg_72_30fab105208816ae;

ARCHITECTURE bmg_72_30fab105208816ae_a OF bmg_72_30fab105208816ae IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_30fab105208816ae
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_30fab105208816ae USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_30fab105208816ae.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 9,
      c_read_width_b => 9,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 9,
      c_write_width_b => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_30fab105208816ae
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_30fab105208816ae_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_8bdf24f02e925a98.vhd when simulating
-- the core, bmg_72_8bdf24f02e925a98. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_8bdf24f02e925a98 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END bmg_72_8bdf24f02e925a98;

ARCHITECTURE bmg_72_8bdf24f02e925a98_a OF bmg_72_8bdf24f02e925a98 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_8bdf24f02e925a98
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_8bdf24f02e925a98 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 3,
      c_addrb_width => 3,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_8bdf24f02e925a98.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 8,
      c_read_depth_b => 8,
      c_read_width_a => 32,
      c_read_width_b => 32,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 8,
      c_write_depth_b => 8,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 32,
      c_write_width_b => 32,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_8bdf24f02e925a98
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_8bdf24f02e925a98_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_d44417b0abe027bf.vhd when simulating
-- the core, bmg_72_d44417b0abe027bf. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_d44417b0abe027bf IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END bmg_72_d44417b0abe027bf;

ARCHITECTURE bmg_72_d44417b0abe027bf_a OF bmg_72_d44417b0abe027bf IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_d44417b0abe027bf
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_d44417b0abe027bf USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_d44417b0abe027bf.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 64,
      c_read_depth_b => 64,
      c_read_width_a => 32,
      c_read_width_b => 32,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 64,
      c_write_depth_b => 64,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 32,
      c_write_width_b => 32,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_d44417b0abe027bf
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_d44417b0abe027bf_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_e4abe4c74ea5aa02.vhd when simulating
-- the core, bmg_72_e4abe4c74ea5aa02. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_e4abe4c74ea5aa02 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END bmg_72_e4abe4c74ea5aa02;

ARCHITECTURE bmg_72_e4abe4c74ea5aa02_a OF bmg_72_e4abe4c74ea5aa02 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_e4abe4c74ea5aa02
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_e4abe4c74ea5aa02 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_e4abe4c74ea5aa02.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 64,
      c_read_depth_b => 64,
      c_read_width_a => 32,
      c_read_width_b => 32,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 64,
      c_write_depth_b => 64,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 32,
      c_write_width_b => 32,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_e4abe4c74ea5aa02
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_e4abe4c74ea5aa02_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_36e2bb554c95560d.vhd when simulating
-- the core, cntr_11_0_36e2bb554c95560d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_36e2bb554c95560d IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END cntr_11_0_36e2bb554c95560d;

ARCHITECTURE cntr_11_0_36e2bb554c95560d_a OF cntr_11_0_36e2bb554c95560d IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_36e2bb554c95560d
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_36e2bb554c95560d USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_36e2bb554c95560d
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_36e2bb554c95560d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_511eb7a1af6f3f2a.vhd when simulating
-- the core, cntr_11_0_511eb7a1af6f3f2a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_511eb7a1af6f3f2a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END cntr_11_0_511eb7a1af6f3f2a;

ARCHITECTURE cntr_11_0_511eb7a1af6f3f2a_a OF cntr_11_0_511eb7a1af6f3f2a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_511eb7a1af6f3f2a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_511eb7a1af6f3f2a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 10,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_511eb7a1af6f3f2a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_511eb7a1af6f3f2a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_6454489cfe866515.vhd when simulating
-- the core, cntr_11_0_6454489cfe866515. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_6454489cfe866515 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END cntr_11_0_6454489cfe866515;

ARCHITECTURE cntr_11_0_6454489cfe866515_a OF cntr_11_0_6454489cfe866515 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_6454489cfe866515
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_6454489cfe866515 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 2,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_6454489cfe866515
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_6454489cfe866515_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_86806e294f737f4c.vhd when simulating
-- the core, cntr_11_0_86806e294f737f4c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_86806e294f737f4c IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_86806e294f737f4c;

ARCHITECTURE cntr_11_0_86806e294f737f4c_a OF cntr_11_0_86806e294f737f4c IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_86806e294f737f4c
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_86806e294f737f4c USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_86806e294f737f4c
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_86806e294f737f4c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_87d991c7bcfe987f.vhd when simulating
-- the core, cntr_11_0_87d991c7bcfe987f. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_87d991c7bcfe987f IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END cntr_11_0_87d991c7bcfe987f;

ARCHITECTURE cntr_11_0_87d991c7bcfe987f_a OF cntr_11_0_87d991c7bcfe987f IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_87d991c7bcfe987f
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_87d991c7bcfe987f USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 5,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_87d991c7bcfe987f
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_87d991c7bcfe987f_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_bcc28bfecf25caff.vhd when simulating
-- the core, cntr_11_0_bcc28bfecf25caff. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_bcc28bfecf25caff IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END cntr_11_0_bcc28bfecf25caff;

ARCHITECTURE cntr_11_0_bcc28bfecf25caff_a OF cntr_11_0_bcc28bfecf25caff IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_bcc28bfecf25caff
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_bcc28bfecf25caff USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 3,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_bcc28bfecf25caff
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_bcc28bfecf25caff_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_d5912692bc2e79ac.vhd when simulating
-- the core, cntr_11_0_d5912692bc2e79ac. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_d5912692bc2e79ac IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
  );
END cntr_11_0_d5912692bc2e79ac;

ARCHITECTURE cntr_11_0_d5912692bc2e79ac_a OF cntr_11_0_d5912692bc2e79ac IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_d5912692bc2e79ac
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_d5912692bc2e79ac USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 15,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_d5912692bc2e79ac
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_d5912692bc2e79ac_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_f068fb73312ae1e5.vhd when simulating
-- the core, cntr_11_0_f068fb73312ae1e5. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_f068fb73312ae1e5 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END cntr_11_0_f068fb73312ae1e5;

ARCHITECTURE cntr_11_0_f068fb73312ae1e5_a OF cntr_11_0_f068fb73312ae1e5 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_f068fb73312ae1e5
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_f068fb73312ae1e5 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 6,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_f068fb73312ae1e5
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_f068fb73312ae1e5_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_06262d82a068201e.vhd when simulating
-- the core, dmg_72_06262d82a068201e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_06262d82a068201e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END dmg_72_06262d82a068201e;

ARCHITECTURE dmg_72_06262d82a068201e_a OF dmg_72_06262d82a068201e IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_06262d82a068201e
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_06262d82a068201e USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 8,
      c_default_data => "0",
      c_depth => 256,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_06262d82a068201e.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 8
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_06262d82a068201e
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_06262d82a068201e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_134e91999cae8947.vhd when simulating
-- the core, dmg_72_134e91999cae8947. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_134e91999cae8947 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END dmg_72_134e91999cae8947;

ARCHITECTURE dmg_72_134e91999cae8947_a OF dmg_72_134e91999cae8947 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_134e91999cae8947
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_134e91999cae8947 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 8,
      c_default_data => "0",
      c_depth => 256,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_134e91999cae8947.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 32
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_134e91999cae8947
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_134e91999cae8947_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_2b0650236539a42c.vhd when simulating
-- the core, dmg_72_2b0650236539a42c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_2b0650236539a42c IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_2b0650236539a42c;

ARCHITECTURE dmg_72_2b0650236539a42c_a OF dmg_72_2b0650236539a42c IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_2b0650236539a42c
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_2b0650236539a42c USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 9,
      c_default_data => "0",
      c_depth => 512,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_2b0650236539a42c.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_2b0650236539a42c
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_2b0650236539a42c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_2be916f69ff4e5b8.vhd when simulating
-- the core, dmg_72_2be916f69ff4e5b8. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_2be916f69ff4e5b8 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_2be916f69ff4e5b8;

ARCHITECTURE dmg_72_2be916f69ff4e5b8_a OF dmg_72_2be916f69ff4e5b8 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_2be916f69ff4e5b8
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_2be916f69ff4e5b8 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 7,
      c_default_data => "0",
      c_depth => 128,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_2be916f69ff4e5b8.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_2be916f69ff4e5b8
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_2be916f69ff4e5b8_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_48a0132db6517610.vhd when simulating
-- the core, dmg_72_48a0132db6517610. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_48a0132db6517610 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_48a0132db6517610;

ARCHITECTURE dmg_72_48a0132db6517610_a OF dmg_72_48a0132db6517610 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_48a0132db6517610
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_48a0132db6517610 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 7,
      c_default_data => "0",
      c_depth => 128,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_48a0132db6517610.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_48a0132db6517610
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_48a0132db6517610_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_58f1077b49388e77.vhd when simulating
-- the core, dmg_72_58f1077b49388e77. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_58f1077b49388e77 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END dmg_72_58f1077b49388e77;

ARCHITECTURE dmg_72_58f1077b49388e77_a OF dmg_72_58f1077b49388e77 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_58f1077b49388e77
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_58f1077b49388e77 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 6,
      c_default_data => "0",
      c_depth => 64,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_58f1077b49388e77.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 7
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_58f1077b49388e77
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_58f1077b49388e77_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_d16d082a6bc00ceb.vhd when simulating
-- the core, dmg_72_d16d082a6bc00ceb. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_d16d082a6bc00ceb IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_d16d082a6bc00ceb;

ARCHITECTURE dmg_72_d16d082a6bc00ceb_a OF dmg_72_d16d082a6bc00ceb IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_d16d082a6bc00ceb
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_d16d082a6bc00ceb USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 9,
      c_default_data => "0",
      c_depth => 512,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_d16d082a6bc00ceb.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_d16d082a6bc00ceb
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_d16d082a6bc00ceb_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_d59da422e431313e.vhd when simulating
-- the core, dmg_72_d59da422e431313e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_d59da422e431313e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END dmg_72_d59da422e431313e;

ARCHITECTURE dmg_72_d59da422e431313e_a OF dmg_72_d59da422e431313e IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_d59da422e431313e
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_d59da422e431313e USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 6,
      c_default_data => "0",
      c_depth => 64,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_d59da422e431313e.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 7
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_d59da422e431313e
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_d59da422e431313e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fifo_fg92_6a1156e8dc43a711.vhd when simulating
-- the core, fifo_fg92_6a1156e8dc43a711. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fifo_fg92_6a1156e8dc43a711 IS
  PORT (
    clk : IN STD_LOGIC;
    srst : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC;
    data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END fifo_fg92_6a1156e8dc43a711;

ARCHITECTURE fifo_fg92_6a1156e8dc43a711_a OF fifo_fg92_6a1156e8dc43a711 IS
-- synthesis translate_off
COMPONENT wrapped_fifo_fg92_6a1156e8dc43a711
  PORT (
    clk : IN STD_LOGIC;
    srst : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC;
    data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fifo_fg92_6a1156e8dc43a711 USE ENTITY XilinxCoreLib.fifo_generator_v9_3(behavioral)
    GENERIC MAP (
      c_add_ngc_constraint => 0,
      c_application_type_axis => 0,
      c_application_type_rach => 0,
      c_application_type_rdch => 0,
      c_application_type_wach => 0,
      c_application_type_wdch => 0,
      c_application_type_wrch => 0,
      c_axi_addr_width => 32,
      c_axi_aruser_width => 1,
      c_axi_awuser_width => 1,
      c_axi_buser_width => 1,
      c_axi_data_width => 64,
      c_axi_id_width => 4,
      c_axi_ruser_width => 1,
      c_axi_type => 0,
      c_axi_wuser_width => 1,
      c_axis_tdata_width => 64,
      c_axis_tdest_width => 4,
      c_axis_tid_width => 8,
      c_axis_tkeep_width => 4,
      c_axis_tstrb_width => 4,
      c_axis_tuser_width => 4,
      c_axis_type => 0,
      c_common_clock => 1,
      c_count_type => 0,
      c_data_count_width => 8,
      c_default_value => "BlankString",
      c_din_width => 32,
      c_din_width_axis => 1,
      c_din_width_rach => 32,
      c_din_width_rdch => 64,
      c_din_width_wach => 32,
      c_din_width_wdch => 64,
      c_din_width_wrch => 2,
      c_dout_rst_val => "0",
      c_dout_width => 32,
      c_enable_rlocs => 0,
      c_enable_rst_sync => 1,
      c_error_injection_type => 0,
      c_error_injection_type_axis => 0,
      c_error_injection_type_rach => 0,
      c_error_injection_type_rdch => 0,
      c_error_injection_type_wach => 0,
      c_error_injection_type_wdch => 0,
      c_error_injection_type_wrch => 0,
      c_family => "virtex6",
      c_full_flags_rst_val => 0,
      c_has_almost_empty => 0,
      c_has_almost_full => 0,
      c_has_axi_aruser => 0,
      c_has_axi_awuser => 0,
      c_has_axi_buser => 0,
      c_has_axi_rd_channel => 0,
      c_has_axi_ruser => 0,
      c_has_axi_wr_channel => 0,
      c_has_axi_wuser => 0,
      c_has_axis_tdata => 0,
      c_has_axis_tdest => 0,
      c_has_axis_tid => 0,
      c_has_axis_tkeep => 0,
      c_has_axis_tlast => 0,
      c_has_axis_tready => 1,
      c_has_axis_tstrb => 0,
      c_has_axis_tuser => 0,
      c_has_backup => 0,
      c_has_data_count => 1,
      c_has_data_counts_axis => 0,
      c_has_data_counts_rach => 0,
      c_has_data_counts_rdch => 0,
      c_has_data_counts_wach => 0,
      c_has_data_counts_wdch => 0,
      c_has_data_counts_wrch => 0,
      c_has_int_clk => 0,
      c_has_master_ce => 0,
      c_has_meminit_file => 0,
      c_has_overflow => 0,
      c_has_prog_flags_axis => 0,
      c_has_prog_flags_rach => 0,
      c_has_prog_flags_rdch => 0,
      c_has_prog_flags_wach => 0,
      c_has_prog_flags_wdch => 0,
      c_has_prog_flags_wrch => 0,
      c_has_rd_data_count => 0,
      c_has_rd_rst => 0,
      c_has_rst => 0,
      c_has_slave_ce => 0,
      c_has_srst => 1,
      c_has_underflow => 0,
      c_has_valid => 0,
      c_has_wr_ack => 0,
      c_has_wr_data_count => 0,
      c_has_wr_rst => 0,
      c_implementation_type => 0,
      c_implementation_type_axis => 1,
      c_implementation_type_rach => 1,
      c_implementation_type_rdch => 1,
      c_implementation_type_wach => 1,
      c_implementation_type_wdch => 1,
      c_implementation_type_wrch => 1,
      c_init_wr_pntr_val => 0,
      c_interface_type => 0,
      c_memory_type => 1,
      c_mif_file_name => "BlankString",
      c_msgon_val => 1,
      c_optimization_mode => 0,
      c_overflow_low => 0,
      c_preload_latency => 2,
      c_preload_regs => 1,
      c_prim_fifo_type => "512x36",
      c_prog_empty_thresh_assert_val => 2,
      c_prog_empty_thresh_assert_val_axis => 1022,
      c_prog_empty_thresh_assert_val_rach => 1022,
      c_prog_empty_thresh_assert_val_rdch => 1022,
      c_prog_empty_thresh_assert_val_wach => 1022,
      c_prog_empty_thresh_assert_val_wdch => 1022,
      c_prog_empty_thresh_assert_val_wrch => 1022,
      c_prog_empty_thresh_negate_val => 3,
      c_prog_empty_type => 0,
      c_prog_empty_type_axis => 0,
      c_prog_empty_type_rach => 0,
      c_prog_empty_type_rdch => 0,
      c_prog_empty_type_wach => 0,
      c_prog_empty_type_wdch => 0,
      c_prog_empty_type_wrch => 0,
      c_prog_full_thresh_assert_val => 254,
      c_prog_full_thresh_assert_val_axis => 1023,
      c_prog_full_thresh_assert_val_rach => 1023,
      c_prog_full_thresh_assert_val_rdch => 1023,
      c_prog_full_thresh_assert_val_wach => 1023,
      c_prog_full_thresh_assert_val_wdch => 1023,
      c_prog_full_thresh_assert_val_wrch => 1023,
      c_prog_full_thresh_negate_val => 253,
      c_prog_full_type => 0,
      c_prog_full_type_axis => 0,
      c_prog_full_type_rach => 0,
      c_prog_full_type_rdch => 0,
      c_prog_full_type_wach => 0,
      c_prog_full_type_wdch => 0,
      c_prog_full_type_wrch => 0,
      c_rach_type => 0,
      c_rd_data_count_width => 8,
      c_rd_depth => 256,
      c_rd_freq => 1,
      c_rd_pntr_width => 8,
      c_rdch_type => 0,
      c_reg_slice_mode_axis => 0,
      c_reg_slice_mode_rach => 0,
      c_reg_slice_mode_rdch => 0,
      c_reg_slice_mode_wach => 0,
      c_reg_slice_mode_wdch => 0,
      c_reg_slice_mode_wrch => 0,
      c_synchronizer_stage => 2,
      c_underflow_low => 0,
      c_use_common_overflow => 0,
      c_use_common_underflow => 0,
      c_use_default_settings => 0,
      c_use_dout_rst => 1,
      c_use_ecc => 0,
      c_use_ecc_axis => 0,
      c_use_ecc_rach => 0,
      c_use_ecc_rdch => 0,
      c_use_ecc_wach => 0,
      c_use_ecc_wdch => 0,
      c_use_ecc_wrch => 0,
      c_use_embedded_reg => 1,
      c_use_fifo16_flags => 0,
      c_use_fwft_data_count => 0,
      c_valid_low => 0,
      c_wach_type => 0,
      c_wdch_type => 0,
      c_wr_ack_low => 0,
      c_wr_data_count_width => 8,
      c_wr_depth => 256,
      c_wr_depth_axis => 1024,
      c_wr_depth_rach => 16,
      c_wr_depth_rdch => 1024,
      c_wr_depth_wach => 16,
      c_wr_depth_wdch => 1024,
      c_wr_depth_wrch => 16,
      c_wr_freq => 1,
      c_wr_pntr_width => 8,
      c_wr_pntr_width_axis => 10,
      c_wr_pntr_width_rach => 4,
      c_wr_pntr_width_rdch => 10,
      c_wr_pntr_width_wach => 4,
      c_wr_pntr_width_wdch => 10,
      c_wr_pntr_width_wrch => 4,
      c_wr_response_latency => 1,
      c_wrch_type => 0
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fifo_fg92_6a1156e8dc43a711
  PORT MAP (
    clk => clk,
    srst => srst,
    din => din,
    wr_en => wr_en,
    rd_en => rd_en,
    dout => dout,
    full => full,
    empty => empty,
    data_count => data_count
  );
-- synthesis translate_on

END fifo_fg92_6a1156e8dc43a711_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_414c0fa5acc33f35.vhd when simulating
-- the core, mult_11_2_414c0fa5acc33f35. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_414c0fa5acc33f35 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END mult_11_2_414c0fa5acc33f35;

ARCHITECTURE mult_11_2_414c0fa5acc33f35_a OF mult_11_2_414c0fa5acc33f35 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_414c0fa5acc33f35
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_414c0fa5acc33f35 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 0,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_zero_detect => 0,
      c_latency => 0,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 31,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_414c0fa5acc33f35
  PORT MAP (
    a => a,
    b => b,
    p => p
  );
-- synthesis translate_on

END mult_11_2_414c0fa5acc33f35_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2015 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_f2bb5a57782af7d9.vhd when simulating
-- the core, mult_11_2_f2bb5a57782af7d9. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_f2bb5a57782af7d9 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END mult_11_2_f2bb5a57782af7d9;

ARCHITECTURE mult_11_2_f2bb5a57782af7d9_a OF mult_11_2_f2bb5a57782af7d9 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_f2bb5a57782af7d9
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_f2bb5a57782af7d9 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 16,
      c_b_type => 1,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_zero_detect => 0,
      c_latency => 0,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 31,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_f2bb5a57782af7d9
  PORT MAP (
    a => a,
    b => b,
    p => p
  );
-- synthesis translate_on

END mult_11_2_f2bb5a57782af7d9_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2012 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: P.49d
--  \   \         Application: netgen
--  /   /         Filename: xfft_v8_0_3683b4047ed128ab.vhd
-- /___/   /\     Timestamp: Wed Jan 27 22:34:22 2016
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -w -sim -ofmt vhdl C:/Users/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c837ea2ae66681b2d/tmp/_cg/xfft_v8_0_3683b4047ed128ab.ngc C:/Users/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c837ea2ae66681b2d/tmp/_cg/xfft_v8_0_3683b4047ed128ab.vhd 
-- Device	: 6vlx240tff1156-2
-- Input file	: C:/Users/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c837ea2ae66681b2d/tmp/_cg/xfft_v8_0_3683b4047ed128ab.ngc
-- Output file	: C:/Users/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c837ea2ae66681b2d/tmp/_cg/xfft_v8_0_3683b4047ed128ab.vhd
-- # of Entities	: 1
-- Design Name	: xfft_v8_0_3683b4047ed128ab
-- Xilinx	: s:\xilinx\14.4\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity xfft_v8_0_3683b4047ed128ab is
  port (
    aclk : in STD_LOGIC := 'X'; 
    aclken : in STD_LOGIC := 'X'; 
    aresetn : in STD_LOGIC := 'X'; 
    s_axis_config_tvalid : in STD_LOGIC := 'X'; 
    s_axis_data_tvalid : in STD_LOGIC := 'X'; 
    s_axis_data_tlast : in STD_LOGIC := 'X'; 
    m_axis_data_tready : in STD_LOGIC := 'X'; 
    m_axis_status_tready : in STD_LOGIC := 'X'; 
    s_axis_config_tready : out STD_LOGIC; 
    s_axis_data_tready : out STD_LOGIC; 
    m_axis_data_tvalid : out STD_LOGIC; 
    m_axis_data_tlast : out STD_LOGIC; 
    m_axis_status_tvalid : out STD_LOGIC; 
    event_frame_started : out STD_LOGIC; 
    event_tlast_unexpected : out STD_LOGIC; 
    event_tlast_missing : out STD_LOGIC; 
    event_fft_overflow : out STD_LOGIC; 
    event_status_channel_halt : out STD_LOGIC; 
    event_data_in_channel_halt : out STD_LOGIC; 
    event_data_out_channel_halt : out STD_LOGIC; 
    s_axis_config_tdata : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    s_axis_data_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    m_axis_data_tdata : out STD_LOGIC_VECTOR ( 31 downto 0 ); 
    m_axis_data_tuser : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    m_axis_status_tdata : out STD_LOGIC_VECTOR ( 7 downto 0 ) 
  );
end xfft_v8_0_3683b4047ed128ab;

architecture STRUCTURE of xfft_v8_0_3683b4047ed128ab is
  signal NlwRenamedSig_OI_m_axis_data_tuser_10_Q : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_data_tuser_8_Q : STD_LOGIC; 
  signal NlwRenamedSig_OI_s_axis_config_tready : STD_LOGIC; 
  signal NlwRenamedSig_OI_s_axis_data_tready : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_data_tvalid : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_status_tvalid : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_frame_started : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_tlast_missing : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_fft_overflow : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_status_channel_halt : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_data_in_channel_halt : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_data_out_channel_halt : STD_LOGIC; 
  signal blk00000001_sig00000fd4 : STD_LOGIC; 
  signal blk00000001_sig00000fd3 : STD_LOGIC; 
  signal blk00000001_sig00000fd2 : STD_LOGIC; 
  signal blk00000001_sig00000fd1 : STD_LOGIC; 
  signal blk00000001_sig00000fd0 : STD_LOGIC; 
  signal blk00000001_sig00000fcf : STD_LOGIC; 
  signal blk00000001_sig00000fce : STD_LOGIC; 
  signal blk00000001_sig00000fcd : STD_LOGIC; 
  signal blk00000001_sig00000fcc : STD_LOGIC; 
  signal blk00000001_sig00000fcb : STD_LOGIC; 
  signal blk00000001_sig00000fca : STD_LOGIC; 
  signal blk00000001_sig00000fc9 : STD_LOGIC; 
  signal blk00000001_sig00000fc8 : STD_LOGIC; 
  signal blk00000001_sig00000fc7 : STD_LOGIC; 
  signal blk00000001_sig00000fc6 : STD_LOGIC; 
  signal blk00000001_sig00000fc5 : STD_LOGIC; 
  signal blk00000001_sig00000fc4 : STD_LOGIC; 
  signal blk00000001_sig00000fc3 : STD_LOGIC; 
  signal blk00000001_sig00000fc2 : STD_LOGIC; 
  signal blk00000001_sig00000fc1 : STD_LOGIC; 
  signal blk00000001_sig00000fc0 : STD_LOGIC; 
  signal blk00000001_sig00000fbf : STD_LOGIC; 
  signal blk00000001_sig00000fbe : STD_LOGIC; 
  signal blk00000001_sig00000fbd : STD_LOGIC; 
  signal blk00000001_sig00000fbc : STD_LOGIC; 
  signal blk00000001_sig00000fbb : STD_LOGIC; 
  signal blk00000001_sig00000fba : STD_LOGIC; 
  signal blk00000001_sig00000fb9 : STD_LOGIC; 
  signal blk00000001_sig00000fb8 : STD_LOGIC; 
  signal blk00000001_sig00000fb7 : STD_LOGIC; 
  signal blk00000001_sig00000fb6 : STD_LOGIC; 
  signal blk00000001_sig00000fb5 : STD_LOGIC; 
  signal blk00000001_sig00000fb4 : STD_LOGIC; 
  signal blk00000001_sig00000fb3 : STD_LOGIC; 
  signal blk00000001_sig00000fb2 : STD_LOGIC; 
  signal blk00000001_sig00000fb1 : STD_LOGIC; 
  signal blk00000001_sig00000fb0 : STD_LOGIC; 
  signal blk00000001_sig00000faf : STD_LOGIC; 
  signal blk00000001_sig00000fae : STD_LOGIC; 
  signal blk00000001_sig00000fad : STD_LOGIC; 
  signal blk00000001_sig00000fac : STD_LOGIC; 
  signal blk00000001_sig00000fab : STD_LOGIC; 
  signal blk00000001_sig00000faa : STD_LOGIC; 
  signal blk00000001_sig00000fa9 : STD_LOGIC; 
  signal blk00000001_sig00000fa8 : STD_LOGIC; 
  signal blk00000001_sig00000fa7 : STD_LOGIC; 
  signal blk00000001_sig00000fa6 : STD_LOGIC; 
  signal blk00000001_sig00000fa5 : STD_LOGIC; 
  signal blk00000001_sig00000fa4 : STD_LOGIC; 
  signal blk00000001_sig00000fa3 : STD_LOGIC; 
  signal blk00000001_sig00000fa2 : STD_LOGIC; 
  signal blk00000001_sig00000fa1 : STD_LOGIC; 
  signal blk00000001_sig00000fa0 : STD_LOGIC; 
  signal blk00000001_sig00000f9f : STD_LOGIC; 
  signal blk00000001_sig00000f9e : STD_LOGIC; 
  signal blk00000001_sig00000f9d : STD_LOGIC; 
  signal blk00000001_sig00000f9c : STD_LOGIC; 
  signal blk00000001_sig00000f9b : STD_LOGIC; 
  signal blk00000001_sig00000f9a : STD_LOGIC; 
  signal blk00000001_sig00000f99 : STD_LOGIC; 
  signal blk00000001_sig00000f98 : STD_LOGIC; 
  signal blk00000001_sig00000f97 : STD_LOGIC; 
  signal blk00000001_sig00000f96 : STD_LOGIC; 
  signal blk00000001_sig00000f95 : STD_LOGIC; 
  signal blk00000001_sig00000f94 : STD_LOGIC; 
  signal blk00000001_sig00000f93 : STD_LOGIC; 
  signal blk00000001_sig00000f92 : STD_LOGIC; 
  signal blk00000001_sig00000f91 : STD_LOGIC; 
  signal blk00000001_sig00000f90 : STD_LOGIC; 
  signal blk00000001_sig00000f8f : STD_LOGIC; 
  signal blk00000001_sig00000f8e : STD_LOGIC; 
  signal blk00000001_sig00000f8d : STD_LOGIC; 
  signal blk00000001_sig00000f8c : STD_LOGIC; 
  signal blk00000001_sig00000f8b : STD_LOGIC; 
  signal blk00000001_sig00000f8a : STD_LOGIC; 
  signal blk00000001_sig00000f89 : STD_LOGIC; 
  signal blk00000001_sig00000f88 : STD_LOGIC; 
  signal blk00000001_sig00000f87 : STD_LOGIC; 
  signal blk00000001_sig00000f86 : STD_LOGIC; 
  signal blk00000001_sig00000f85 : STD_LOGIC; 
  signal blk00000001_sig00000f84 : STD_LOGIC; 
  signal blk00000001_sig00000f83 : STD_LOGIC; 
  signal blk00000001_sig00000f82 : STD_LOGIC; 
  signal blk00000001_sig00000f81 : STD_LOGIC; 
  signal blk00000001_sig00000f80 : STD_LOGIC; 
  signal blk00000001_sig00000f7f : STD_LOGIC; 
  signal blk00000001_sig00000f7e : STD_LOGIC; 
  signal blk00000001_sig00000f7d : STD_LOGIC; 
  signal blk00000001_sig00000f7c : STD_LOGIC; 
  signal blk00000001_sig00000f7b : STD_LOGIC; 
  signal blk00000001_sig00000f7a : STD_LOGIC; 
  signal blk00000001_sig00000f79 : STD_LOGIC; 
  signal blk00000001_sig00000f78 : STD_LOGIC; 
  signal blk00000001_sig00000f77 : STD_LOGIC; 
  signal blk00000001_sig00000f76 : STD_LOGIC; 
  signal blk00000001_sig00000f75 : STD_LOGIC; 
  signal blk00000001_sig00000f74 : STD_LOGIC; 
  signal blk00000001_sig00000f73 : STD_LOGIC; 
  signal blk00000001_sig00000f72 : STD_LOGIC; 
  signal blk00000001_sig00000f71 : STD_LOGIC; 
  signal blk00000001_sig00000f70 : STD_LOGIC; 
  signal blk00000001_sig00000f6f : STD_LOGIC; 
  signal blk00000001_sig00000f6e : STD_LOGIC; 
  signal blk00000001_sig00000f6d : STD_LOGIC; 
  signal blk00000001_sig00000f6c : STD_LOGIC; 
  signal blk00000001_sig00000f6b : STD_LOGIC; 
  signal blk00000001_sig00000f6a : STD_LOGIC; 
  signal blk00000001_sig00000f69 : STD_LOGIC; 
  signal blk00000001_sig00000f68 : STD_LOGIC; 
  signal blk00000001_sig00000f67 : STD_LOGIC; 
  signal blk00000001_sig00000f66 : STD_LOGIC; 
  signal blk00000001_sig00000f65 : STD_LOGIC; 
  signal blk00000001_sig00000f64 : STD_LOGIC; 
  signal blk00000001_sig00000f63 : STD_LOGIC; 
  signal blk00000001_sig00000f62 : STD_LOGIC; 
  signal blk00000001_sig00000f61 : STD_LOGIC; 
  signal blk00000001_sig00000f60 : STD_LOGIC; 
  signal blk00000001_sig00000f5f : STD_LOGIC; 
  signal blk00000001_sig00000f5e : STD_LOGIC; 
  signal blk00000001_sig00000f5d : STD_LOGIC; 
  signal blk00000001_sig00000f5c : STD_LOGIC; 
  signal blk00000001_sig00000f5b : STD_LOGIC; 
  signal blk00000001_sig00000f5a : STD_LOGIC; 
  signal blk00000001_sig00000f59 : STD_LOGIC; 
  signal blk00000001_sig00000f58 : STD_LOGIC; 
  signal blk00000001_sig00000f57 : STD_LOGIC; 
  signal blk00000001_sig00000f56 : STD_LOGIC; 
  signal blk00000001_sig00000f55 : STD_LOGIC; 
  signal blk00000001_sig00000f54 : STD_LOGIC; 
  signal blk00000001_sig00000f53 : STD_LOGIC; 
  signal blk00000001_sig00000f52 : STD_LOGIC; 
  signal blk00000001_sig00000f51 : STD_LOGIC; 
  signal blk00000001_sig00000f50 : STD_LOGIC; 
  signal blk00000001_sig00000f4f : STD_LOGIC; 
  signal blk00000001_sig00000f4e : STD_LOGIC; 
  signal blk00000001_sig00000f4d : STD_LOGIC; 
  signal blk00000001_sig00000f4c : STD_LOGIC; 
  signal blk00000001_sig00000f4b : STD_LOGIC; 
  signal blk00000001_sig00000f4a : STD_LOGIC; 
  signal blk00000001_sig00000f49 : STD_LOGIC; 
  signal blk00000001_sig00000f48 : STD_LOGIC; 
  signal blk00000001_sig00000f47 : STD_LOGIC; 
  signal blk00000001_sig00000f46 : STD_LOGIC; 
  signal blk00000001_sig00000f45 : STD_LOGIC; 
  signal blk00000001_sig00000f44 : STD_LOGIC; 
  signal blk00000001_sig00000f43 : STD_LOGIC; 
  signal blk00000001_sig00000f42 : STD_LOGIC; 
  signal blk00000001_sig00000f41 : STD_LOGIC; 
  signal blk00000001_sig00000f40 : STD_LOGIC; 
  signal blk00000001_sig00000f3f : STD_LOGIC; 
  signal blk00000001_sig00000f3e : STD_LOGIC; 
  signal blk00000001_sig00000f3d : STD_LOGIC; 
  signal blk00000001_sig00000f3c : STD_LOGIC; 
  signal blk00000001_sig00000f3b : STD_LOGIC; 
  signal blk00000001_sig00000f3a : STD_LOGIC; 
  signal blk00000001_sig00000f39 : STD_LOGIC; 
  signal blk00000001_sig00000f38 : STD_LOGIC; 
  signal blk00000001_sig00000f37 : STD_LOGIC; 
  signal blk00000001_sig00000f36 : STD_LOGIC; 
  signal blk00000001_sig00000f35 : STD_LOGIC; 
  signal blk00000001_sig00000f34 : STD_LOGIC; 
  signal blk00000001_sig00000f33 : STD_LOGIC; 
  signal blk00000001_sig00000f32 : STD_LOGIC; 
  signal blk00000001_sig00000f31 : STD_LOGIC; 
  signal blk00000001_sig00000f30 : STD_LOGIC; 
  signal blk00000001_sig00000f2f : STD_LOGIC; 
  signal blk00000001_sig00000f2e : STD_LOGIC; 
  signal blk00000001_sig00000f2d : STD_LOGIC; 
  signal blk00000001_sig00000f2c : STD_LOGIC; 
  signal blk00000001_sig00000f2b : STD_LOGIC; 
  signal blk00000001_sig00000f2a : STD_LOGIC; 
  signal blk00000001_sig00000f29 : STD_LOGIC; 
  signal blk00000001_sig00000f28 : STD_LOGIC; 
  signal blk00000001_sig00000f27 : STD_LOGIC; 
  signal blk00000001_sig00000f26 : STD_LOGIC; 
  signal blk00000001_sig00000f25 : STD_LOGIC; 
  signal blk00000001_sig00000f24 : STD_LOGIC; 
  signal blk00000001_sig00000f23 : STD_LOGIC; 
  signal blk00000001_sig00000f22 : STD_LOGIC; 
  signal blk00000001_sig00000f21 : STD_LOGIC; 
  signal blk00000001_sig00000f20 : STD_LOGIC; 
  signal blk00000001_sig00000f1f : STD_LOGIC; 
  signal blk00000001_sig00000f1e : STD_LOGIC; 
  signal blk00000001_sig00000f1d : STD_LOGIC; 
  signal blk00000001_sig00000f1c : STD_LOGIC; 
  signal blk00000001_sig00000f1b : STD_LOGIC; 
  signal blk00000001_sig00000f1a : STD_LOGIC; 
  signal blk00000001_sig00000f19 : STD_LOGIC; 
  signal blk00000001_sig00000f18 : STD_LOGIC; 
  signal blk00000001_sig00000f17 : STD_LOGIC; 
  signal blk00000001_sig00000f16 : STD_LOGIC; 
  signal blk00000001_sig00000f15 : STD_LOGIC; 
  signal blk00000001_sig00000f14 : STD_LOGIC; 
  signal blk00000001_sig00000f13 : STD_LOGIC; 
  signal blk00000001_sig00000f12 : STD_LOGIC; 
  signal blk00000001_sig00000f11 : STD_LOGIC; 
  signal blk00000001_sig00000f10 : STD_LOGIC; 
  signal blk00000001_sig00000f0f : STD_LOGIC; 
  signal blk00000001_sig00000f0e : STD_LOGIC; 
  signal blk00000001_sig00000f0d : STD_LOGIC; 
  signal blk00000001_sig00000f0c : STD_LOGIC; 
  signal blk00000001_sig00000f0b : STD_LOGIC; 
  signal blk00000001_sig00000f0a : STD_LOGIC; 
  signal blk00000001_sig00000f09 : STD_LOGIC; 
  signal blk00000001_sig00000f08 : STD_LOGIC; 
  signal blk00000001_sig00000f07 : STD_LOGIC; 
  signal blk00000001_sig00000f06 : STD_LOGIC; 
  signal blk00000001_sig00000f05 : STD_LOGIC; 
  signal blk00000001_sig00000f04 : STD_LOGIC; 
  signal blk00000001_sig00000f03 : STD_LOGIC; 
  signal blk00000001_sig00000f02 : STD_LOGIC; 
  signal blk00000001_sig00000f01 : STD_LOGIC; 
  signal blk00000001_sig00000f00 : STD_LOGIC; 
  signal blk00000001_sig00000eff : STD_LOGIC; 
  signal blk00000001_sig00000efe : STD_LOGIC; 
  signal blk00000001_sig00000efd : STD_LOGIC; 
  signal blk00000001_sig00000efc : STD_LOGIC; 
  signal blk00000001_sig00000efb : STD_LOGIC; 
  signal blk00000001_sig00000efa : STD_LOGIC; 
  signal blk00000001_sig00000ef9 : STD_LOGIC; 
  signal blk00000001_sig00000ef8 : STD_LOGIC; 
  signal blk00000001_sig00000ef7 : STD_LOGIC; 
  signal blk00000001_sig00000ef6 : STD_LOGIC; 
  signal blk00000001_sig00000ef5 : STD_LOGIC; 
  signal blk00000001_sig00000ef4 : STD_LOGIC; 
  signal blk00000001_sig00000ef3 : STD_LOGIC; 
  signal blk00000001_sig00000ef2 : STD_LOGIC; 
  signal blk00000001_sig00000ef1 : STD_LOGIC; 
  signal blk00000001_sig00000ef0 : STD_LOGIC; 
  signal blk00000001_sig00000eef : STD_LOGIC; 
  signal blk00000001_sig00000eee : STD_LOGIC; 
  signal blk00000001_sig00000eed : STD_LOGIC; 
  signal blk00000001_sig00000eec : STD_LOGIC; 
  signal blk00000001_sig00000eeb : STD_LOGIC; 
  signal blk00000001_sig00000eea : STD_LOGIC; 
  signal blk00000001_sig00000ee9 : STD_LOGIC; 
  signal blk00000001_sig00000ee8 : STD_LOGIC; 
  signal blk00000001_sig00000ee7 : STD_LOGIC; 
  signal blk00000001_sig00000ee6 : STD_LOGIC; 
  signal blk00000001_sig00000ee5 : STD_LOGIC; 
  signal blk00000001_sig00000ee4 : STD_LOGIC; 
  signal blk00000001_sig00000ee3 : STD_LOGIC; 
  signal blk00000001_sig00000ee2 : STD_LOGIC; 
  signal blk00000001_sig00000ee1 : STD_LOGIC; 
  signal blk00000001_sig00000ee0 : STD_LOGIC; 
  signal blk00000001_sig00000edf : STD_LOGIC; 
  signal blk00000001_sig00000ede : STD_LOGIC; 
  signal blk00000001_sig00000edd : STD_LOGIC; 
  signal blk00000001_sig00000edc : STD_LOGIC; 
  signal blk00000001_sig00000edb : STD_LOGIC; 
  signal blk00000001_sig00000eda : STD_LOGIC; 
  signal blk00000001_sig00000ed9 : STD_LOGIC; 
  signal blk00000001_sig00000ed8 : STD_LOGIC; 
  signal blk00000001_sig00000ed7 : STD_LOGIC; 
  signal blk00000001_sig00000ed6 : STD_LOGIC; 
  signal blk00000001_sig00000ed5 : STD_LOGIC; 
  signal blk00000001_sig00000ed4 : STD_LOGIC; 
  signal blk00000001_sig00000ed3 : STD_LOGIC; 
  signal blk00000001_sig00000ed2 : STD_LOGIC; 
  signal blk00000001_sig00000ed1 : STD_LOGIC; 
  signal blk00000001_sig00000ed0 : STD_LOGIC; 
  signal blk00000001_sig00000ecf : STD_LOGIC; 
  signal blk00000001_sig00000ece : STD_LOGIC; 
  signal blk00000001_sig00000ecd : STD_LOGIC; 
  signal blk00000001_sig00000ecc : STD_LOGIC; 
  signal blk00000001_sig00000ecb : STD_LOGIC; 
  signal blk00000001_sig00000eca : STD_LOGIC; 
  signal blk00000001_sig00000ec9 : STD_LOGIC; 
  signal blk00000001_sig00000ec8 : STD_LOGIC; 
  signal blk00000001_sig00000ec7 : STD_LOGIC; 
  signal blk00000001_sig00000ec6 : STD_LOGIC; 
  signal blk00000001_sig00000ec5 : STD_LOGIC; 
  signal blk00000001_sig00000ec4 : STD_LOGIC; 
  signal blk00000001_sig00000ec3 : STD_LOGIC; 
  signal blk00000001_sig00000ec2 : STD_LOGIC; 
  signal blk00000001_sig00000ec1 : STD_LOGIC; 
  signal blk00000001_sig00000ec0 : STD_LOGIC; 
  signal blk00000001_sig00000ebf : STD_LOGIC; 
  signal blk00000001_sig00000ebe : STD_LOGIC; 
  signal blk00000001_sig00000ebd : STD_LOGIC; 
  signal blk00000001_sig00000ebc : STD_LOGIC; 
  signal blk00000001_sig00000ebb : STD_LOGIC; 
  signal blk00000001_sig00000eba : STD_LOGIC; 
  signal blk00000001_sig00000eb9 : STD_LOGIC; 
  signal blk00000001_sig00000eb8 : STD_LOGIC; 
  signal blk00000001_sig00000eb7 : STD_LOGIC; 
  signal blk00000001_sig00000eb6 : STD_LOGIC; 
  signal blk00000001_sig00000eb5 : STD_LOGIC; 
  signal blk00000001_sig00000eb4 : STD_LOGIC; 
  signal blk00000001_sig00000eb3 : STD_LOGIC; 
  signal blk00000001_sig00000eb2 : STD_LOGIC; 
  signal blk00000001_sig00000eb1 : STD_LOGIC; 
  signal blk00000001_sig00000eb0 : STD_LOGIC; 
  signal blk00000001_sig00000eaf : STD_LOGIC; 
  signal blk00000001_sig00000eae : STD_LOGIC; 
  signal blk00000001_sig00000ead : STD_LOGIC; 
  signal blk00000001_sig00000eac : STD_LOGIC; 
  signal blk00000001_sig00000eab : STD_LOGIC; 
  signal blk00000001_sig00000eaa : STD_LOGIC; 
  signal blk00000001_sig00000ea9 : STD_LOGIC; 
  signal blk00000001_sig00000ea8 : STD_LOGIC; 
  signal blk00000001_sig00000ea7 : STD_LOGIC; 
  signal blk00000001_sig00000ea6 : STD_LOGIC; 
  signal blk00000001_sig00000ea5 : STD_LOGIC; 
  signal blk00000001_sig00000ea4 : STD_LOGIC; 
  signal blk00000001_sig00000ea3 : STD_LOGIC; 
  signal blk00000001_sig00000ea2 : STD_LOGIC; 
  signal blk00000001_sig00000ea1 : STD_LOGIC; 
  signal blk00000001_sig00000ea0 : STD_LOGIC; 
  signal blk00000001_sig00000e9f : STD_LOGIC; 
  signal blk00000001_sig00000e9e : STD_LOGIC; 
  signal blk00000001_sig00000e9d : STD_LOGIC; 
  signal blk00000001_sig00000e9c : STD_LOGIC; 
  signal blk00000001_sig00000e9b : STD_LOGIC; 
  signal blk00000001_sig00000e9a : STD_LOGIC; 
  signal blk00000001_sig00000e99 : STD_LOGIC; 
  signal blk00000001_sig00000e98 : STD_LOGIC; 
  signal blk00000001_sig00000e97 : STD_LOGIC; 
  signal blk00000001_sig00000e96 : STD_LOGIC; 
  signal blk00000001_sig00000e95 : STD_LOGIC; 
  signal blk00000001_sig00000e94 : STD_LOGIC; 
  signal blk00000001_sig00000e93 : STD_LOGIC; 
  signal blk00000001_sig00000e92 : STD_LOGIC; 
  signal blk00000001_sig00000e91 : STD_LOGIC; 
  signal blk00000001_sig00000e90 : STD_LOGIC; 
  signal blk00000001_sig00000e8f : STD_LOGIC; 
  signal blk00000001_sig00000e8e : STD_LOGIC; 
  signal blk00000001_sig00000e8d : STD_LOGIC; 
  signal blk00000001_sig00000e8c : STD_LOGIC; 
  signal blk00000001_sig00000e8b : STD_LOGIC; 
  signal blk00000001_sig00000e8a : STD_LOGIC; 
  signal blk00000001_sig00000e89 : STD_LOGIC; 
  signal blk00000001_sig00000e88 : STD_LOGIC; 
  signal blk00000001_sig00000e87 : STD_LOGIC; 
  signal blk00000001_sig00000e86 : STD_LOGIC; 
  signal blk00000001_sig00000e85 : STD_LOGIC; 
  signal blk00000001_sig00000e84 : STD_LOGIC; 
  signal blk00000001_sig00000e83 : STD_LOGIC; 
  signal blk00000001_sig00000e82 : STD_LOGIC; 
  signal blk00000001_sig00000e81 : STD_LOGIC; 
  signal blk00000001_sig00000e80 : STD_LOGIC; 
  signal blk00000001_sig00000e7f : STD_LOGIC; 
  signal blk00000001_sig00000e7e : STD_LOGIC; 
  signal blk00000001_sig00000e7d : STD_LOGIC; 
  signal blk00000001_sig00000e7c : STD_LOGIC; 
  signal blk00000001_sig00000e7b : STD_LOGIC; 
  signal blk00000001_sig00000e7a : STD_LOGIC; 
  signal blk00000001_sig00000e79 : STD_LOGIC; 
  signal blk00000001_sig00000e78 : STD_LOGIC; 
  signal blk00000001_sig00000e77 : STD_LOGIC; 
  signal blk00000001_sig00000e76 : STD_LOGIC; 
  signal blk00000001_sig00000e75 : STD_LOGIC; 
  signal blk00000001_sig00000e74 : STD_LOGIC; 
  signal blk00000001_sig00000e73 : STD_LOGIC; 
  signal blk00000001_sig00000e72 : STD_LOGIC; 
  signal blk00000001_sig00000e71 : STD_LOGIC; 
  signal blk00000001_sig00000e70 : STD_LOGIC; 
  signal blk00000001_sig00000e6f : STD_LOGIC; 
  signal blk00000001_sig00000e6e : STD_LOGIC; 
  signal blk00000001_sig00000e6d : STD_LOGIC; 
  signal blk00000001_sig00000e6c : STD_LOGIC; 
  signal blk00000001_sig00000e6b : STD_LOGIC; 
  signal blk00000001_sig00000e6a : STD_LOGIC; 
  signal blk00000001_sig00000e69 : STD_LOGIC; 
  signal blk00000001_sig00000e68 : STD_LOGIC; 
  signal blk00000001_sig00000e67 : STD_LOGIC; 
  signal blk00000001_sig00000e66 : STD_LOGIC; 
  signal blk00000001_sig00000e65 : STD_LOGIC; 
  signal blk00000001_sig00000e64 : STD_LOGIC; 
  signal blk00000001_sig00000e63 : STD_LOGIC; 
  signal blk00000001_sig00000e62 : STD_LOGIC; 
  signal blk00000001_sig00000e61 : STD_LOGIC; 
  signal blk00000001_sig00000e60 : STD_LOGIC; 
  signal blk00000001_sig00000e5f : STD_LOGIC; 
  signal blk00000001_sig00000e5e : STD_LOGIC; 
  signal blk00000001_sig00000e5d : STD_LOGIC; 
  signal blk00000001_sig00000e5c : STD_LOGIC; 
  signal blk00000001_sig00000e5b : STD_LOGIC; 
  signal blk00000001_sig00000e5a : STD_LOGIC; 
  signal blk00000001_sig00000e59 : STD_LOGIC; 
  signal blk00000001_sig00000e58 : STD_LOGIC; 
  signal blk00000001_sig00000e57 : STD_LOGIC; 
  signal blk00000001_sig00000e56 : STD_LOGIC; 
  signal blk00000001_sig00000e55 : STD_LOGIC; 
  signal blk00000001_sig00000e54 : STD_LOGIC; 
  signal blk00000001_sig00000e53 : STD_LOGIC; 
  signal blk00000001_sig00000e52 : STD_LOGIC; 
  signal blk00000001_sig00000e51 : STD_LOGIC; 
  signal blk00000001_sig00000e50 : STD_LOGIC; 
  signal blk00000001_sig00000e4f : STD_LOGIC; 
  signal blk00000001_sig00000e4e : STD_LOGIC; 
  signal blk00000001_sig00000e4d : STD_LOGIC; 
  signal blk00000001_sig00000e4c : STD_LOGIC; 
  signal blk00000001_sig00000e4b : STD_LOGIC; 
  signal blk00000001_sig00000e4a : STD_LOGIC; 
  signal blk00000001_sig00000e49 : STD_LOGIC; 
  signal blk00000001_sig00000e48 : STD_LOGIC; 
  signal blk00000001_sig00000e47 : STD_LOGIC; 
  signal blk00000001_sig00000e46 : STD_LOGIC; 
  signal blk00000001_sig00000e45 : STD_LOGIC; 
  signal blk00000001_sig00000e44 : STD_LOGIC; 
  signal blk00000001_sig00000e43 : STD_LOGIC; 
  signal blk00000001_sig00000e42 : STD_LOGIC; 
  signal blk00000001_sig00000e41 : STD_LOGIC; 
  signal blk00000001_sig00000e40 : STD_LOGIC; 
  signal blk00000001_sig00000e3f : STD_LOGIC; 
  signal blk00000001_sig00000e3e : STD_LOGIC; 
  signal blk00000001_sig00000e3d : STD_LOGIC; 
  signal blk00000001_sig00000e3c : STD_LOGIC; 
  signal blk00000001_sig00000e3b : STD_LOGIC; 
  signal blk00000001_sig00000e3a : STD_LOGIC; 
  signal blk00000001_sig00000e39 : STD_LOGIC; 
  signal blk00000001_sig00000e38 : STD_LOGIC; 
  signal blk00000001_sig00000e37 : STD_LOGIC; 
  signal blk00000001_sig00000e36 : STD_LOGIC; 
  signal blk00000001_sig00000e35 : STD_LOGIC; 
  signal blk00000001_sig00000e34 : STD_LOGIC; 
  signal blk00000001_sig00000e33 : STD_LOGIC; 
  signal blk00000001_sig00000e32 : STD_LOGIC; 
  signal blk00000001_sig00000e31 : STD_LOGIC; 
  signal blk00000001_sig00000e30 : STD_LOGIC; 
  signal blk00000001_sig00000e2f : STD_LOGIC; 
  signal blk00000001_sig00000e2e : STD_LOGIC; 
  signal blk00000001_sig00000e2d : STD_LOGIC; 
  signal blk00000001_sig00000e2c : STD_LOGIC; 
  signal blk00000001_sig00000e2b : STD_LOGIC; 
  signal blk00000001_sig00000e2a : STD_LOGIC; 
  signal blk00000001_sig00000e29 : STD_LOGIC; 
  signal blk00000001_sig00000e28 : STD_LOGIC; 
  signal blk00000001_sig00000e27 : STD_LOGIC; 
  signal blk00000001_sig00000e26 : STD_LOGIC; 
  signal blk00000001_sig00000e25 : STD_LOGIC; 
  signal blk00000001_sig00000e24 : STD_LOGIC; 
  signal blk00000001_sig00000e23 : STD_LOGIC; 
  signal blk00000001_sig00000e22 : STD_LOGIC; 
  signal blk00000001_sig00000e21 : STD_LOGIC; 
  signal blk00000001_sig00000e20 : STD_LOGIC; 
  signal blk00000001_sig00000e1f : STD_LOGIC; 
  signal blk00000001_sig00000e1e : STD_LOGIC; 
  signal blk00000001_sig00000e1d : STD_LOGIC; 
  signal blk00000001_sig00000e1c : STD_LOGIC; 
  signal blk00000001_sig00000e1b : STD_LOGIC; 
  signal blk00000001_sig00000e1a : STD_LOGIC; 
  signal blk00000001_sig00000e19 : STD_LOGIC; 
  signal blk00000001_sig00000e18 : STD_LOGIC; 
  signal blk00000001_sig00000e17 : STD_LOGIC; 
  signal blk00000001_sig00000e16 : STD_LOGIC; 
  signal blk00000001_sig00000e15 : STD_LOGIC; 
  signal blk00000001_sig00000e14 : STD_LOGIC; 
  signal blk00000001_sig00000e13 : STD_LOGIC; 
  signal blk00000001_sig00000e12 : STD_LOGIC; 
  signal blk00000001_sig00000e11 : STD_LOGIC; 
  signal blk00000001_sig00000e10 : STD_LOGIC; 
  signal blk00000001_sig00000e0f : STD_LOGIC; 
  signal blk00000001_sig00000e0e : STD_LOGIC; 
  signal blk00000001_sig00000e0d : STD_LOGIC; 
  signal blk00000001_sig00000e0c : STD_LOGIC; 
  signal blk00000001_sig00000e0b : STD_LOGIC; 
  signal blk00000001_sig00000e0a : STD_LOGIC; 
  signal blk00000001_sig00000e09 : STD_LOGIC; 
  signal blk00000001_sig00000e08 : STD_LOGIC; 
  signal blk00000001_sig00000e07 : STD_LOGIC; 
  signal blk00000001_sig00000e06 : STD_LOGIC; 
  signal blk00000001_sig00000e05 : STD_LOGIC; 
  signal blk00000001_sig00000e04 : STD_LOGIC; 
  signal blk00000001_sig00000e03 : STD_LOGIC; 
  signal blk00000001_sig00000e02 : STD_LOGIC; 
  signal blk00000001_sig00000e01 : STD_LOGIC; 
  signal blk00000001_sig00000e00 : STD_LOGIC; 
  signal blk00000001_sig00000dff : STD_LOGIC; 
  signal blk00000001_sig00000dfe : STD_LOGIC; 
  signal blk00000001_sig00000dfd : STD_LOGIC; 
  signal blk00000001_sig00000dfc : STD_LOGIC; 
  signal blk00000001_sig00000dfb : STD_LOGIC; 
  signal blk00000001_sig00000dfa : STD_LOGIC; 
  signal blk00000001_sig00000df9 : STD_LOGIC; 
  signal blk00000001_sig00000df8 : STD_LOGIC; 
  signal blk00000001_sig00000df7 : STD_LOGIC; 
  signal blk00000001_sig00000df6 : STD_LOGIC; 
  signal blk00000001_sig00000df5 : STD_LOGIC; 
  signal blk00000001_sig00000df4 : STD_LOGIC; 
  signal blk00000001_sig00000df3 : STD_LOGIC; 
  signal blk00000001_sig00000df2 : STD_LOGIC; 
  signal blk00000001_sig00000df1 : STD_LOGIC; 
  signal blk00000001_sig00000df0 : STD_LOGIC; 
  signal blk00000001_sig00000def : STD_LOGIC; 
  signal blk00000001_sig00000dee : STD_LOGIC; 
  signal blk00000001_sig00000ded : STD_LOGIC; 
  signal blk00000001_sig00000dec : STD_LOGIC; 
  signal blk00000001_sig00000deb : STD_LOGIC; 
  signal blk00000001_sig00000dea : STD_LOGIC; 
  signal blk00000001_sig00000de9 : STD_LOGIC; 
  signal blk00000001_sig00000de8 : STD_LOGIC; 
  signal blk00000001_sig00000de7 : STD_LOGIC; 
  signal blk00000001_sig00000de6 : STD_LOGIC; 
  signal blk00000001_sig00000de5 : STD_LOGIC; 
  signal blk00000001_sig00000de4 : STD_LOGIC; 
  signal blk00000001_sig00000de3 : STD_LOGIC; 
  signal blk00000001_sig00000de2 : STD_LOGIC; 
  signal blk00000001_sig00000de1 : STD_LOGIC; 
  signal blk00000001_sig00000de0 : STD_LOGIC; 
  signal blk00000001_sig00000ddf : STD_LOGIC; 
  signal blk00000001_sig00000dde : STD_LOGIC; 
  signal blk00000001_sig00000ddd : STD_LOGIC; 
  signal blk00000001_sig00000ddc : STD_LOGIC; 
  signal blk00000001_sig00000ddb : STD_LOGIC; 
  signal blk00000001_sig00000dda : STD_LOGIC; 
  signal blk00000001_sig00000dd9 : STD_LOGIC; 
  signal blk00000001_sig00000dd8 : STD_LOGIC; 
  signal blk00000001_sig00000dd7 : STD_LOGIC; 
  signal blk00000001_sig00000dd6 : STD_LOGIC; 
  signal blk00000001_sig00000dd5 : STD_LOGIC; 
  signal blk00000001_sig00000dd4 : STD_LOGIC; 
  signal blk00000001_sig00000dd3 : STD_LOGIC; 
  signal blk00000001_sig00000dd2 : STD_LOGIC; 
  signal blk00000001_sig00000dd1 : STD_LOGIC; 
  signal blk00000001_sig00000dd0 : STD_LOGIC; 
  signal blk00000001_sig00000dcf : STD_LOGIC; 
  signal blk00000001_sig00000dce : STD_LOGIC; 
  signal blk00000001_sig00000dcd : STD_LOGIC; 
  signal blk00000001_sig00000dcc : STD_LOGIC; 
  signal blk00000001_sig00000dcb : STD_LOGIC; 
  signal blk00000001_sig00000dca : STD_LOGIC; 
  signal blk00000001_sig00000dc9 : STD_LOGIC; 
  signal blk00000001_sig00000dc8 : STD_LOGIC; 
  signal blk00000001_sig00000dc7 : STD_LOGIC; 
  signal blk00000001_sig00000dc6 : STD_LOGIC; 
  signal blk00000001_sig00000dc5 : STD_LOGIC; 
  signal blk00000001_sig00000dc4 : STD_LOGIC; 
  signal blk00000001_sig00000dc3 : STD_LOGIC; 
  signal blk00000001_sig00000dc2 : STD_LOGIC; 
  signal blk00000001_sig00000dc1 : STD_LOGIC; 
  signal blk00000001_sig00000dc0 : STD_LOGIC; 
  signal blk00000001_sig00000dbf : STD_LOGIC; 
  signal blk00000001_sig00000dbe : STD_LOGIC; 
  signal blk00000001_sig00000dbd : STD_LOGIC; 
  signal blk00000001_sig00000dbc : STD_LOGIC; 
  signal blk00000001_sig00000dbb : STD_LOGIC; 
  signal blk00000001_sig00000dba : STD_LOGIC; 
  signal blk00000001_sig00000db9 : STD_LOGIC; 
  signal blk00000001_sig00000db8 : STD_LOGIC; 
  signal blk00000001_sig00000db7 : STD_LOGIC; 
  signal blk00000001_sig00000db6 : STD_LOGIC; 
  signal blk00000001_sig00000db5 : STD_LOGIC; 
  signal blk00000001_sig00000db4 : STD_LOGIC; 
  signal blk00000001_sig00000db3 : STD_LOGIC; 
  signal blk00000001_sig00000db2 : STD_LOGIC; 
  signal blk00000001_sig00000db1 : STD_LOGIC; 
  signal blk00000001_sig00000db0 : STD_LOGIC; 
  signal blk00000001_sig00000daf : STD_LOGIC; 
  signal blk00000001_sig00000dae : STD_LOGIC; 
  signal blk00000001_sig00000dad : STD_LOGIC; 
  signal blk00000001_sig00000dac : STD_LOGIC; 
  signal blk00000001_sig00000dab : STD_LOGIC; 
  signal blk00000001_sig00000daa : STD_LOGIC; 
  signal blk00000001_sig00000da9 : STD_LOGIC; 
  signal blk00000001_sig00000da8 : STD_LOGIC; 
  signal blk00000001_sig00000da7 : STD_LOGIC; 
  signal blk00000001_sig00000da6 : STD_LOGIC; 
  signal blk00000001_sig00000da5 : STD_LOGIC; 
  signal blk00000001_sig00000da4 : STD_LOGIC; 
  signal blk00000001_sig00000da3 : STD_LOGIC; 
  signal blk00000001_sig00000da2 : STD_LOGIC; 
  signal blk00000001_sig00000da1 : STD_LOGIC; 
  signal blk00000001_sig00000da0 : STD_LOGIC; 
  signal blk00000001_sig00000d9f : STD_LOGIC; 
  signal blk00000001_sig00000d9e : STD_LOGIC; 
  signal blk00000001_sig00000d9d : STD_LOGIC; 
  signal blk00000001_sig00000d9c : STD_LOGIC; 
  signal blk00000001_sig00000d9b : STD_LOGIC; 
  signal blk00000001_sig00000d9a : STD_LOGIC; 
  signal blk00000001_sig00000d99 : STD_LOGIC; 
  signal blk00000001_sig00000d98 : STD_LOGIC; 
  signal blk00000001_sig00000d97 : STD_LOGIC; 
  signal blk00000001_sig00000d96 : STD_LOGIC; 
  signal blk00000001_sig00000d95 : STD_LOGIC; 
  signal blk00000001_sig00000d94 : STD_LOGIC; 
  signal blk00000001_sig00000d93 : STD_LOGIC; 
  signal blk00000001_sig00000d92 : STD_LOGIC; 
  signal blk00000001_sig00000d91 : STD_LOGIC; 
  signal blk00000001_sig00000d90 : STD_LOGIC; 
  signal blk00000001_sig00000d8f : STD_LOGIC; 
  signal blk00000001_sig00000d8e : STD_LOGIC; 
  signal blk00000001_sig00000d8d : STD_LOGIC; 
  signal blk00000001_sig00000d8c : STD_LOGIC; 
  signal blk00000001_sig00000d8b : STD_LOGIC; 
  signal blk00000001_sig00000d8a : STD_LOGIC; 
  signal blk00000001_sig00000d89 : STD_LOGIC; 
  signal blk00000001_sig00000d88 : STD_LOGIC; 
  signal blk00000001_sig00000d87 : STD_LOGIC; 
  signal blk00000001_sig00000d86 : STD_LOGIC; 
  signal blk00000001_sig00000d85 : STD_LOGIC; 
  signal blk00000001_sig00000d84 : STD_LOGIC; 
  signal blk00000001_sig00000d83 : STD_LOGIC; 
  signal blk00000001_sig00000d82 : STD_LOGIC; 
  signal blk00000001_sig00000d81 : STD_LOGIC; 
  signal blk00000001_sig00000d80 : STD_LOGIC; 
  signal blk00000001_sig00000d7f : STD_LOGIC; 
  signal blk00000001_sig00000d7e : STD_LOGIC; 
  signal blk00000001_sig00000d7d : STD_LOGIC; 
  signal blk00000001_sig00000d7c : STD_LOGIC; 
  signal blk00000001_sig00000d7b : STD_LOGIC; 
  signal blk00000001_sig00000d7a : STD_LOGIC; 
  signal blk00000001_sig00000d79 : STD_LOGIC; 
  signal blk00000001_sig00000d78 : STD_LOGIC; 
  signal blk00000001_sig00000d77 : STD_LOGIC; 
  signal blk00000001_sig00000d76 : STD_LOGIC; 
  signal blk00000001_sig00000d75 : STD_LOGIC; 
  signal blk00000001_sig00000d74 : STD_LOGIC; 
  signal blk00000001_sig00000d73 : STD_LOGIC; 
  signal blk00000001_sig00000d72 : STD_LOGIC; 
  signal blk00000001_sig00000d71 : STD_LOGIC; 
  signal blk00000001_sig00000d70 : STD_LOGIC; 
  signal blk00000001_sig00000d6f : STD_LOGIC; 
  signal blk00000001_sig00000d6e : STD_LOGIC; 
  signal blk00000001_sig00000d6d : STD_LOGIC; 
  signal blk00000001_sig00000d6c : STD_LOGIC; 
  signal blk00000001_sig00000d6b : STD_LOGIC; 
  signal blk00000001_sig00000d6a : STD_LOGIC; 
  signal blk00000001_sig00000d69 : STD_LOGIC; 
  signal blk00000001_sig00000d68 : STD_LOGIC; 
  signal blk00000001_sig00000d67 : STD_LOGIC; 
  signal blk00000001_sig00000d66 : STD_LOGIC; 
  signal blk00000001_sig00000d65 : STD_LOGIC; 
  signal blk00000001_sig00000d64 : STD_LOGIC; 
  signal blk00000001_sig00000d63 : STD_LOGIC; 
  signal blk00000001_sig00000d62 : STD_LOGIC; 
  signal blk00000001_sig00000d61 : STD_LOGIC; 
  signal blk00000001_sig00000d60 : STD_LOGIC; 
  signal blk00000001_sig00000d5f : STD_LOGIC; 
  signal blk00000001_sig00000d5e : STD_LOGIC; 
  signal blk00000001_sig00000d5d : STD_LOGIC; 
  signal blk00000001_sig00000d5c : STD_LOGIC; 
  signal blk00000001_sig00000d5b : STD_LOGIC; 
  signal blk00000001_sig00000d5a : STD_LOGIC; 
  signal blk00000001_sig00000d59 : STD_LOGIC; 
  signal blk00000001_sig00000d58 : STD_LOGIC; 
  signal blk00000001_sig00000d57 : STD_LOGIC; 
  signal blk00000001_sig00000d56 : STD_LOGIC; 
  signal blk00000001_sig00000d55 : STD_LOGIC; 
  signal blk00000001_sig00000d54 : STD_LOGIC; 
  signal blk00000001_sig00000d53 : STD_LOGIC; 
  signal blk00000001_sig00000d52 : STD_LOGIC; 
  signal blk00000001_sig00000d51 : STD_LOGIC; 
  signal blk00000001_sig00000d50 : STD_LOGIC; 
  signal blk00000001_sig00000d4f : STD_LOGIC; 
  signal blk00000001_sig00000d4e : STD_LOGIC; 
  signal blk00000001_sig00000d4d : STD_LOGIC; 
  signal blk00000001_sig00000d4c : STD_LOGIC; 
  signal blk00000001_sig00000d4b : STD_LOGIC; 
  signal blk00000001_sig00000d4a : STD_LOGIC; 
  signal blk00000001_sig00000d49 : STD_LOGIC; 
  signal blk00000001_sig00000d48 : STD_LOGIC; 
  signal blk00000001_sig00000d47 : STD_LOGIC; 
  signal blk00000001_sig00000d46 : STD_LOGIC; 
  signal blk00000001_sig00000d45 : STD_LOGIC; 
  signal blk00000001_sig00000d44 : STD_LOGIC; 
  signal blk00000001_sig00000d43 : STD_LOGIC; 
  signal blk00000001_sig00000d42 : STD_LOGIC; 
  signal blk00000001_sig00000d41 : STD_LOGIC; 
  signal blk00000001_sig00000d40 : STD_LOGIC; 
  signal blk00000001_sig00000d3f : STD_LOGIC; 
  signal blk00000001_sig00000d3e : STD_LOGIC; 
  signal blk00000001_sig00000d3d : STD_LOGIC; 
  signal blk00000001_sig00000d3c : STD_LOGIC; 
  signal blk00000001_sig00000d3b : STD_LOGIC; 
  signal blk00000001_sig00000d3a : STD_LOGIC; 
  signal blk00000001_sig00000d39 : STD_LOGIC; 
  signal blk00000001_sig00000d38 : STD_LOGIC; 
  signal blk00000001_sig00000d37 : STD_LOGIC; 
  signal blk00000001_sig00000d36 : STD_LOGIC; 
  signal blk00000001_sig00000d35 : STD_LOGIC; 
  signal blk00000001_sig00000d34 : STD_LOGIC; 
  signal blk00000001_sig00000d33 : STD_LOGIC; 
  signal blk00000001_sig00000d32 : STD_LOGIC; 
  signal blk00000001_sig00000d31 : STD_LOGIC; 
  signal blk00000001_sig00000d30 : STD_LOGIC; 
  signal blk00000001_sig00000d2f : STD_LOGIC; 
  signal blk00000001_sig00000d2e : STD_LOGIC; 
  signal blk00000001_sig00000d2d : STD_LOGIC; 
  signal blk00000001_sig00000d2c : STD_LOGIC; 
  signal blk00000001_sig00000d2b : STD_LOGIC; 
  signal blk00000001_sig00000d2a : STD_LOGIC; 
  signal blk00000001_sig00000d29 : STD_LOGIC; 
  signal blk00000001_sig00000d28 : STD_LOGIC; 
  signal blk00000001_sig00000d27 : STD_LOGIC; 
  signal blk00000001_sig00000d26 : STD_LOGIC; 
  signal blk00000001_sig00000d25 : STD_LOGIC; 
  signal blk00000001_sig00000d24 : STD_LOGIC; 
  signal blk00000001_sig00000d23 : STD_LOGIC; 
  signal blk00000001_sig00000d22 : STD_LOGIC; 
  signal blk00000001_sig00000d21 : STD_LOGIC; 
  signal blk00000001_sig00000d20 : STD_LOGIC; 
  signal blk00000001_sig00000d1f : STD_LOGIC; 
  signal blk00000001_sig00000d1e : STD_LOGIC; 
  signal blk00000001_sig00000d1d : STD_LOGIC; 
  signal blk00000001_sig00000d1c : STD_LOGIC; 
  signal blk00000001_sig00000d1b : STD_LOGIC; 
  signal blk00000001_sig00000d1a : STD_LOGIC; 
  signal blk00000001_sig00000d19 : STD_LOGIC; 
  signal blk00000001_sig00000d18 : STD_LOGIC; 
  signal blk00000001_sig00000d17 : STD_LOGIC; 
  signal blk00000001_sig00000d16 : STD_LOGIC; 
  signal blk00000001_sig00000d15 : STD_LOGIC; 
  signal blk00000001_sig00000d14 : STD_LOGIC; 
  signal blk00000001_sig00000d13 : STD_LOGIC; 
  signal blk00000001_sig00000d12 : STD_LOGIC; 
  signal blk00000001_sig00000d11 : STD_LOGIC; 
  signal blk00000001_sig00000d10 : STD_LOGIC; 
  signal blk00000001_sig00000d0f : STD_LOGIC; 
  signal blk00000001_sig00000d0e : STD_LOGIC; 
  signal blk00000001_sig00000d0d : STD_LOGIC; 
  signal blk00000001_sig00000d0c : STD_LOGIC; 
  signal blk00000001_sig00000d0b : STD_LOGIC; 
  signal blk00000001_sig00000d0a : STD_LOGIC; 
  signal blk00000001_sig00000d09 : STD_LOGIC; 
  signal blk00000001_sig00000d08 : STD_LOGIC; 
  signal blk00000001_sig00000d07 : STD_LOGIC; 
  signal blk00000001_sig00000d06 : STD_LOGIC; 
  signal blk00000001_sig00000d05 : STD_LOGIC; 
  signal blk00000001_sig00000d04 : STD_LOGIC; 
  signal blk00000001_sig00000d03 : STD_LOGIC; 
  signal blk00000001_sig00000d02 : STD_LOGIC; 
  signal blk00000001_sig00000d01 : STD_LOGIC; 
  signal blk00000001_sig00000d00 : STD_LOGIC; 
  signal blk00000001_sig00000cff : STD_LOGIC; 
  signal blk00000001_sig00000cfe : STD_LOGIC; 
  signal blk00000001_sig00000cfd : STD_LOGIC; 
  signal blk00000001_sig00000cfc : STD_LOGIC; 
  signal blk00000001_sig00000cfb : STD_LOGIC; 
  signal blk00000001_sig00000cfa : STD_LOGIC; 
  signal blk00000001_sig00000cf9 : STD_LOGIC; 
  signal blk00000001_sig00000cf8 : STD_LOGIC; 
  signal blk00000001_sig00000cf7 : STD_LOGIC; 
  signal blk00000001_sig00000cf6 : STD_LOGIC; 
  signal blk00000001_sig00000cf5 : STD_LOGIC; 
  signal blk00000001_sig00000cf4 : STD_LOGIC; 
  signal blk00000001_sig00000cf3 : STD_LOGIC; 
  signal blk00000001_sig00000cf2 : STD_LOGIC; 
  signal blk00000001_sig00000cf1 : STD_LOGIC; 
  signal blk00000001_sig00000cf0 : STD_LOGIC; 
  signal blk00000001_sig00000cef : STD_LOGIC; 
  signal blk00000001_sig00000cee : STD_LOGIC; 
  signal blk00000001_sig00000ced : STD_LOGIC; 
  signal blk00000001_sig00000cec : STD_LOGIC; 
  signal blk00000001_sig00000ceb : STD_LOGIC; 
  signal blk00000001_sig00000cea : STD_LOGIC; 
  signal blk00000001_sig00000ce9 : STD_LOGIC; 
  signal blk00000001_sig00000ce8 : STD_LOGIC; 
  signal blk00000001_sig00000ce7 : STD_LOGIC; 
  signal blk00000001_sig00000ce6 : STD_LOGIC; 
  signal blk00000001_sig00000ce5 : STD_LOGIC; 
  signal blk00000001_sig00000ce4 : STD_LOGIC; 
  signal blk00000001_sig00000ce3 : STD_LOGIC; 
  signal blk00000001_sig00000ce2 : STD_LOGIC; 
  signal blk00000001_sig00000ce1 : STD_LOGIC; 
  signal blk00000001_sig00000ce0 : STD_LOGIC; 
  signal blk00000001_sig00000cdf : STD_LOGIC; 
  signal blk00000001_sig00000cde : STD_LOGIC; 
  signal blk00000001_sig00000cdd : STD_LOGIC; 
  signal blk00000001_sig00000cdc : STD_LOGIC; 
  signal blk00000001_sig00000cdb : STD_LOGIC; 
  signal blk00000001_sig00000cda : STD_LOGIC; 
  signal blk00000001_sig00000cd9 : STD_LOGIC; 
  signal blk00000001_sig00000cd8 : STD_LOGIC; 
  signal blk00000001_sig00000cd7 : STD_LOGIC; 
  signal blk00000001_sig00000cd6 : STD_LOGIC; 
  signal blk00000001_sig00000cd5 : STD_LOGIC; 
  signal blk00000001_sig00000cd4 : STD_LOGIC; 
  signal blk00000001_sig00000cd3 : STD_LOGIC; 
  signal blk00000001_sig00000cd2 : STD_LOGIC; 
  signal blk00000001_sig00000cd1 : STD_LOGIC; 
  signal blk00000001_sig00000cd0 : STD_LOGIC; 
  signal blk00000001_sig00000ccf : STD_LOGIC; 
  signal blk00000001_sig00000cce : STD_LOGIC; 
  signal blk00000001_sig00000ccd : STD_LOGIC; 
  signal blk00000001_sig00000ccc : STD_LOGIC; 
  signal blk00000001_sig00000ccb : STD_LOGIC; 
  signal blk00000001_sig00000cca : STD_LOGIC; 
  signal blk00000001_sig00000cc9 : STD_LOGIC; 
  signal blk00000001_sig00000cc8 : STD_LOGIC; 
  signal blk00000001_sig00000cc7 : STD_LOGIC; 
  signal blk00000001_sig00000cc6 : STD_LOGIC; 
  signal blk00000001_sig00000cc5 : STD_LOGIC; 
  signal blk00000001_sig00000cc4 : STD_LOGIC; 
  signal blk00000001_sig00000cc3 : STD_LOGIC; 
  signal blk00000001_sig00000cc2 : STD_LOGIC; 
  signal blk00000001_sig00000cc1 : STD_LOGIC; 
  signal blk00000001_sig00000cc0 : STD_LOGIC; 
  signal blk00000001_sig00000cbf : STD_LOGIC; 
  signal blk00000001_sig00000cbe : STD_LOGIC; 
  signal blk00000001_sig00000cbd : STD_LOGIC; 
  signal blk00000001_sig00000cbc : STD_LOGIC; 
  signal blk00000001_sig00000cbb : STD_LOGIC; 
  signal blk00000001_sig00000cba : STD_LOGIC; 
  signal blk00000001_sig00000cb9 : STD_LOGIC; 
  signal blk00000001_sig00000cb8 : STD_LOGIC; 
  signal blk00000001_sig00000cb7 : STD_LOGIC; 
  signal blk00000001_sig00000cb6 : STD_LOGIC; 
  signal blk00000001_sig00000cb5 : STD_LOGIC; 
  signal blk00000001_sig00000cb4 : STD_LOGIC; 
  signal blk00000001_sig00000cb3 : STD_LOGIC; 
  signal blk00000001_sig00000cb2 : STD_LOGIC; 
  signal blk00000001_sig00000cb1 : STD_LOGIC; 
  signal blk00000001_sig00000cb0 : STD_LOGIC; 
  signal blk00000001_sig00000caf : STD_LOGIC; 
  signal blk00000001_sig00000cae : STD_LOGIC; 
  signal blk00000001_sig00000cad : STD_LOGIC; 
  signal blk00000001_sig00000cac : STD_LOGIC; 
  signal blk00000001_sig00000cab : STD_LOGIC; 
  signal blk00000001_sig00000caa : STD_LOGIC; 
  signal blk00000001_sig00000ca9 : STD_LOGIC; 
  signal blk00000001_sig00000ca8 : STD_LOGIC; 
  signal blk00000001_sig00000ca7 : STD_LOGIC; 
  signal blk00000001_sig00000ca6 : STD_LOGIC; 
  signal blk00000001_sig00000ca5 : STD_LOGIC; 
  signal blk00000001_sig00000ca4 : STD_LOGIC; 
  signal blk00000001_sig00000ca3 : STD_LOGIC; 
  signal blk00000001_sig00000ca2 : STD_LOGIC; 
  signal blk00000001_sig00000ca1 : STD_LOGIC; 
  signal blk00000001_sig00000ca0 : STD_LOGIC; 
  signal blk00000001_sig00000c9f : STD_LOGIC; 
  signal blk00000001_sig00000c9e : STD_LOGIC; 
  signal blk00000001_sig00000c9d : STD_LOGIC; 
  signal blk00000001_sig00000c9c : STD_LOGIC; 
  signal blk00000001_sig00000c9b : STD_LOGIC; 
  signal blk00000001_sig00000c9a : STD_LOGIC; 
  signal blk00000001_sig00000c99 : STD_LOGIC; 
  signal blk00000001_sig00000c98 : STD_LOGIC; 
  signal blk00000001_sig00000c97 : STD_LOGIC; 
  signal blk00000001_sig00000c96 : STD_LOGIC; 
  signal blk00000001_sig00000c95 : STD_LOGIC; 
  signal blk00000001_sig00000c94 : STD_LOGIC; 
  signal blk00000001_sig00000c93 : STD_LOGIC; 
  signal blk00000001_sig00000c92 : STD_LOGIC; 
  signal blk00000001_sig00000c91 : STD_LOGIC; 
  signal blk00000001_sig00000c90 : STD_LOGIC; 
  signal blk00000001_sig00000c8f : STD_LOGIC; 
  signal blk00000001_sig00000c8e : STD_LOGIC; 
  signal blk00000001_sig00000c8d : STD_LOGIC; 
  signal blk00000001_sig00000c8c : STD_LOGIC; 
  signal blk00000001_sig00000c8b : STD_LOGIC; 
  signal blk00000001_sig00000c8a : STD_LOGIC; 
  signal blk00000001_sig00000c89 : STD_LOGIC; 
  signal blk00000001_sig00000c88 : STD_LOGIC; 
  signal blk00000001_sig00000c87 : STD_LOGIC; 
  signal blk00000001_sig00000c86 : STD_LOGIC; 
  signal blk00000001_sig00000c85 : STD_LOGIC; 
  signal blk00000001_sig00000c84 : STD_LOGIC; 
  signal blk00000001_sig00000c83 : STD_LOGIC; 
  signal blk00000001_sig00000c82 : STD_LOGIC; 
  signal blk00000001_sig00000c81 : STD_LOGIC; 
  signal blk00000001_sig00000c80 : STD_LOGIC; 
  signal blk00000001_sig00000c7f : STD_LOGIC; 
  signal blk00000001_sig00000c7e : STD_LOGIC; 
  signal blk00000001_sig00000c7d : STD_LOGIC; 
  signal blk00000001_sig00000c7c : STD_LOGIC; 
  signal blk00000001_sig00000c7b : STD_LOGIC; 
  signal blk00000001_sig00000c7a : STD_LOGIC; 
  signal blk00000001_sig00000c79 : STD_LOGIC; 
  signal blk00000001_sig00000c78 : STD_LOGIC; 
  signal blk00000001_sig00000c77 : STD_LOGIC; 
  signal blk00000001_sig00000c76 : STD_LOGIC; 
  signal blk00000001_sig00000c75 : STD_LOGIC; 
  signal blk00000001_sig00000c74 : STD_LOGIC; 
  signal blk00000001_sig00000c73 : STD_LOGIC; 
  signal blk00000001_sig00000c72 : STD_LOGIC; 
  signal blk00000001_sig00000c71 : STD_LOGIC; 
  signal blk00000001_sig00000c70 : STD_LOGIC; 
  signal blk00000001_sig00000c6f : STD_LOGIC; 
  signal blk00000001_sig00000c6e : STD_LOGIC; 
  signal blk00000001_sig00000c6d : STD_LOGIC; 
  signal blk00000001_sig00000c6c : STD_LOGIC; 
  signal blk00000001_sig00000c6b : STD_LOGIC; 
  signal blk00000001_sig00000c6a : STD_LOGIC; 
  signal blk00000001_sig00000c69 : STD_LOGIC; 
  signal blk00000001_sig00000c68 : STD_LOGIC; 
  signal blk00000001_sig00000c67 : STD_LOGIC; 
  signal blk00000001_sig00000c66 : STD_LOGIC; 
  signal blk00000001_sig00000c65 : STD_LOGIC; 
  signal blk00000001_sig00000c64 : STD_LOGIC; 
  signal blk00000001_sig00000c63 : STD_LOGIC; 
  signal blk00000001_sig00000c62 : STD_LOGIC; 
  signal blk00000001_sig00000c61 : STD_LOGIC; 
  signal blk00000001_sig00000c60 : STD_LOGIC; 
  signal blk00000001_sig00000c5f : STD_LOGIC; 
  signal blk00000001_sig00000c5e : STD_LOGIC; 
  signal blk00000001_sig00000c5d : STD_LOGIC; 
  signal blk00000001_sig00000c5c : STD_LOGIC; 
  signal blk00000001_sig00000c5b : STD_LOGIC; 
  signal blk00000001_sig00000c5a : STD_LOGIC; 
  signal blk00000001_sig00000c59 : STD_LOGIC; 
  signal blk00000001_sig00000c58 : STD_LOGIC; 
  signal blk00000001_sig00000c57 : STD_LOGIC; 
  signal blk00000001_sig00000c56 : STD_LOGIC; 
  signal blk00000001_sig00000c55 : STD_LOGIC; 
  signal blk00000001_sig00000c54 : STD_LOGIC; 
  signal blk00000001_sig00000c53 : STD_LOGIC; 
  signal blk00000001_sig00000c52 : STD_LOGIC; 
  signal blk00000001_sig00000c51 : STD_LOGIC; 
  signal blk00000001_sig00000c50 : STD_LOGIC; 
  signal blk00000001_sig00000c4f : STD_LOGIC; 
  signal blk00000001_sig00000c4e : STD_LOGIC; 
  signal blk00000001_sig00000c4d : STD_LOGIC; 
  signal blk00000001_sig00000c4c : STD_LOGIC; 
  signal blk00000001_sig00000c4b : STD_LOGIC; 
  signal blk00000001_sig00000c4a : STD_LOGIC; 
  signal blk00000001_sig00000c49 : STD_LOGIC; 
  signal blk00000001_sig00000c48 : STD_LOGIC; 
  signal blk00000001_sig00000c47 : STD_LOGIC; 
  signal blk00000001_sig00000c46 : STD_LOGIC; 
  signal blk00000001_sig00000c45 : STD_LOGIC; 
  signal blk00000001_sig00000c44 : STD_LOGIC; 
  signal blk00000001_sig00000c43 : STD_LOGIC; 
  signal blk00000001_sig00000c42 : STD_LOGIC; 
  signal blk00000001_sig00000c41 : STD_LOGIC; 
  signal blk00000001_sig00000c40 : STD_LOGIC; 
  signal blk00000001_sig00000c3f : STD_LOGIC; 
  signal blk00000001_sig00000c3e : STD_LOGIC; 
  signal blk00000001_sig00000c3d : STD_LOGIC; 
  signal blk00000001_sig00000c3c : STD_LOGIC; 
  signal blk00000001_sig00000c3b : STD_LOGIC; 
  signal blk00000001_sig00000c3a : STD_LOGIC; 
  signal blk00000001_sig00000c39 : STD_LOGIC; 
  signal blk00000001_sig00000c38 : STD_LOGIC; 
  signal blk00000001_sig00000c37 : STD_LOGIC; 
  signal blk00000001_sig00000c36 : STD_LOGIC; 
  signal blk00000001_sig00000c35 : STD_LOGIC; 
  signal blk00000001_sig00000c34 : STD_LOGIC; 
  signal blk00000001_sig00000c33 : STD_LOGIC; 
  signal blk00000001_sig00000c32 : STD_LOGIC; 
  signal blk00000001_sig00000c31 : STD_LOGIC; 
  signal blk00000001_sig00000c30 : STD_LOGIC; 
  signal blk00000001_sig00000c2f : STD_LOGIC; 
  signal blk00000001_sig00000c2e : STD_LOGIC; 
  signal blk00000001_sig00000c2d : STD_LOGIC; 
  signal blk00000001_sig00000c2c : STD_LOGIC; 
  signal blk00000001_sig00000c2b : STD_LOGIC; 
  signal blk00000001_sig00000c2a : STD_LOGIC; 
  signal blk00000001_sig00000c29 : STD_LOGIC; 
  signal blk00000001_sig00000c28 : STD_LOGIC; 
  signal blk00000001_sig00000c27 : STD_LOGIC; 
  signal blk00000001_sig00000c26 : STD_LOGIC; 
  signal blk00000001_sig00000c25 : STD_LOGIC; 
  signal blk00000001_sig00000c24 : STD_LOGIC; 
  signal blk00000001_sig00000c23 : STD_LOGIC; 
  signal blk00000001_sig00000c22 : STD_LOGIC; 
  signal blk00000001_sig00000c21 : STD_LOGIC; 
  signal blk00000001_sig00000c20 : STD_LOGIC; 
  signal blk00000001_sig00000c1f : STD_LOGIC; 
  signal blk00000001_sig00000c1e : STD_LOGIC; 
  signal blk00000001_sig00000c1d : STD_LOGIC; 
  signal blk00000001_sig00000c1c : STD_LOGIC; 
  signal blk00000001_sig00000c1b : STD_LOGIC; 
  signal blk00000001_sig00000c1a : STD_LOGIC; 
  signal blk00000001_sig00000c19 : STD_LOGIC; 
  signal blk00000001_sig00000c18 : STD_LOGIC; 
  signal blk00000001_sig00000c17 : STD_LOGIC; 
  signal blk00000001_sig00000c16 : STD_LOGIC; 
  signal blk00000001_sig00000c15 : STD_LOGIC; 
  signal blk00000001_sig00000c14 : STD_LOGIC; 
  signal blk00000001_sig00000c13 : STD_LOGIC; 
  signal blk00000001_sig00000c12 : STD_LOGIC; 
  signal blk00000001_sig00000c11 : STD_LOGIC; 
  signal blk00000001_sig00000c10 : STD_LOGIC; 
  signal blk00000001_sig00000c0f : STD_LOGIC; 
  signal blk00000001_sig00000c0e : STD_LOGIC; 
  signal blk00000001_sig00000c0d : STD_LOGIC; 
  signal blk00000001_sig00000c0c : STD_LOGIC; 
  signal blk00000001_sig00000c0b : STD_LOGIC; 
  signal blk00000001_sig00000c0a : STD_LOGIC; 
  signal blk00000001_sig00000c09 : STD_LOGIC; 
  signal blk00000001_sig00000c08 : STD_LOGIC; 
  signal blk00000001_sig00000c07 : STD_LOGIC; 
  signal blk00000001_sig00000c06 : STD_LOGIC; 
  signal blk00000001_sig00000c05 : STD_LOGIC; 
  signal blk00000001_sig00000c04 : STD_LOGIC; 
  signal blk00000001_sig00000c03 : STD_LOGIC; 
  signal blk00000001_sig00000c02 : STD_LOGIC; 
  signal blk00000001_sig00000c01 : STD_LOGIC; 
  signal blk00000001_sig00000c00 : STD_LOGIC; 
  signal blk00000001_sig00000bff : STD_LOGIC; 
  signal blk00000001_sig00000bfe : STD_LOGIC; 
  signal blk00000001_sig00000bfd : STD_LOGIC; 
  signal blk00000001_sig00000bfc : STD_LOGIC; 
  signal blk00000001_sig00000bfb : STD_LOGIC; 
  signal blk00000001_sig00000bfa : STD_LOGIC; 
  signal blk00000001_sig00000bf9 : STD_LOGIC; 
  signal blk00000001_sig00000bf8 : STD_LOGIC; 
  signal blk00000001_sig00000bf7 : STD_LOGIC; 
  signal blk00000001_sig00000bf6 : STD_LOGIC; 
  signal blk00000001_sig00000bf5 : STD_LOGIC; 
  signal blk00000001_sig00000bf4 : STD_LOGIC; 
  signal blk00000001_sig00000bf3 : STD_LOGIC; 
  signal blk00000001_sig00000bf2 : STD_LOGIC; 
  signal blk00000001_sig00000bf1 : STD_LOGIC; 
  signal blk00000001_sig00000bf0 : STD_LOGIC; 
  signal blk00000001_sig00000bef : STD_LOGIC; 
  signal blk00000001_sig00000bee : STD_LOGIC; 
  signal blk00000001_sig00000bed : STD_LOGIC; 
  signal blk00000001_sig00000bec : STD_LOGIC; 
  signal blk00000001_sig00000beb : STD_LOGIC; 
  signal blk00000001_sig00000bea : STD_LOGIC; 
  signal blk00000001_sig00000be9 : STD_LOGIC; 
  signal blk00000001_sig00000be8 : STD_LOGIC; 
  signal blk00000001_sig00000be7 : STD_LOGIC; 
  signal blk00000001_sig00000be6 : STD_LOGIC; 
  signal blk00000001_sig00000be5 : STD_LOGIC; 
  signal blk00000001_sig00000be4 : STD_LOGIC; 
  signal blk00000001_sig00000be3 : STD_LOGIC; 
  signal blk00000001_sig00000be2 : STD_LOGIC; 
  signal blk00000001_sig00000be1 : STD_LOGIC; 
  signal blk00000001_sig00000be0 : STD_LOGIC; 
  signal blk00000001_sig00000bdf : STD_LOGIC; 
  signal blk00000001_sig00000bde : STD_LOGIC; 
  signal blk00000001_sig00000bdd : STD_LOGIC; 
  signal blk00000001_sig00000bdc : STD_LOGIC; 
  signal blk00000001_sig00000bdb : STD_LOGIC; 
  signal blk00000001_sig00000bda : STD_LOGIC; 
  signal blk00000001_sig00000bd9 : STD_LOGIC; 
  signal blk00000001_sig00000bd8 : STD_LOGIC; 
  signal blk00000001_sig00000bd7 : STD_LOGIC; 
  signal blk00000001_sig00000bd6 : STD_LOGIC; 
  signal blk00000001_sig00000bd5 : STD_LOGIC; 
  signal blk00000001_sig00000bd4 : STD_LOGIC; 
  signal blk00000001_sig00000bd3 : STD_LOGIC; 
  signal blk00000001_sig00000bd2 : STD_LOGIC; 
  signal blk00000001_sig00000bd1 : STD_LOGIC; 
  signal blk00000001_sig00000bd0 : STD_LOGIC; 
  signal blk00000001_sig00000bcf : STD_LOGIC; 
  signal blk00000001_sig00000bce : STD_LOGIC; 
  signal blk00000001_sig00000bcd : STD_LOGIC; 
  signal blk00000001_sig00000bcc : STD_LOGIC; 
  signal blk00000001_sig00000bcb : STD_LOGIC; 
  signal blk00000001_sig00000bca : STD_LOGIC; 
  signal blk00000001_sig00000bc9 : STD_LOGIC; 
  signal blk00000001_sig00000bc8 : STD_LOGIC; 
  signal blk00000001_sig00000bc7 : STD_LOGIC; 
  signal blk00000001_sig00000bc6 : STD_LOGIC; 
  signal blk00000001_sig00000bc5 : STD_LOGIC; 
  signal blk00000001_sig00000bc4 : STD_LOGIC; 
  signal blk00000001_sig00000bc3 : STD_LOGIC; 
  signal blk00000001_sig00000bc2 : STD_LOGIC; 
  signal blk00000001_sig00000bc1 : STD_LOGIC; 
  signal blk00000001_sig00000bc0 : STD_LOGIC; 
  signal blk00000001_sig00000bbf : STD_LOGIC; 
  signal blk00000001_sig00000bbe : STD_LOGIC; 
  signal blk00000001_sig00000bbd : STD_LOGIC; 
  signal blk00000001_sig00000bbc : STD_LOGIC; 
  signal blk00000001_sig00000bbb : STD_LOGIC; 
  signal blk00000001_sig00000bba : STD_LOGIC; 
  signal blk00000001_sig00000bb9 : STD_LOGIC; 
  signal blk00000001_sig00000bb8 : STD_LOGIC; 
  signal blk00000001_sig00000bb7 : STD_LOGIC; 
  signal blk00000001_sig00000bb6 : STD_LOGIC; 
  signal blk00000001_sig00000bb5 : STD_LOGIC; 
  signal blk00000001_sig00000bb4 : STD_LOGIC; 
  signal blk00000001_sig00000bb3 : STD_LOGIC; 
  signal blk00000001_sig00000bb2 : STD_LOGIC; 
  signal blk00000001_sig00000bb1 : STD_LOGIC; 
  signal blk00000001_sig00000bb0 : STD_LOGIC; 
  signal blk00000001_sig00000baf : STD_LOGIC; 
  signal blk00000001_sig00000bae : STD_LOGIC; 
  signal blk00000001_sig00000bad : STD_LOGIC; 
  signal blk00000001_sig00000bac : STD_LOGIC; 
  signal blk00000001_sig00000bab : STD_LOGIC; 
  signal blk00000001_sig00000baa : STD_LOGIC; 
  signal blk00000001_sig00000ba9 : STD_LOGIC; 
  signal blk00000001_sig00000ba8 : STD_LOGIC; 
  signal blk00000001_sig00000ba7 : STD_LOGIC; 
  signal blk00000001_sig00000ba6 : STD_LOGIC; 
  signal blk00000001_sig00000ba5 : STD_LOGIC; 
  signal blk00000001_sig00000ba4 : STD_LOGIC; 
  signal blk00000001_sig00000ba3 : STD_LOGIC; 
  signal blk00000001_sig00000ba2 : STD_LOGIC; 
  signal blk00000001_sig00000ba1 : STD_LOGIC; 
  signal blk00000001_sig00000ba0 : STD_LOGIC; 
  signal blk00000001_sig00000b9f : STD_LOGIC; 
  signal blk00000001_sig00000b9e : STD_LOGIC; 
  signal blk00000001_sig00000b9d : STD_LOGIC; 
  signal blk00000001_sig00000b9c : STD_LOGIC; 
  signal blk00000001_sig00000b9b : STD_LOGIC; 
  signal blk00000001_sig00000b9a : STD_LOGIC; 
  signal blk00000001_sig00000b99 : STD_LOGIC; 
  signal blk00000001_sig00000b98 : STD_LOGIC; 
  signal blk00000001_sig00000b97 : STD_LOGIC; 
  signal blk00000001_sig00000b96 : STD_LOGIC; 
  signal blk00000001_sig00000b95 : STD_LOGIC; 
  signal blk00000001_sig00000b94 : STD_LOGIC; 
  signal blk00000001_sig00000b93 : STD_LOGIC; 
  signal blk00000001_sig00000b92 : STD_LOGIC; 
  signal blk00000001_sig00000b91 : STD_LOGIC; 
  signal blk00000001_sig00000b90 : STD_LOGIC; 
  signal blk00000001_sig00000b8f : STD_LOGIC; 
  signal blk00000001_sig00000b8e : STD_LOGIC; 
  signal blk00000001_sig00000b8d : STD_LOGIC; 
  signal blk00000001_sig00000b8c : STD_LOGIC; 
  signal blk00000001_sig00000b8b : STD_LOGIC; 
  signal blk00000001_sig00000b8a : STD_LOGIC; 
  signal blk00000001_sig00000b89 : STD_LOGIC; 
  signal blk00000001_sig00000b88 : STD_LOGIC; 
  signal blk00000001_sig00000b87 : STD_LOGIC; 
  signal blk00000001_sig00000b86 : STD_LOGIC; 
  signal blk00000001_sig00000b85 : STD_LOGIC; 
  signal blk00000001_sig00000b84 : STD_LOGIC; 
  signal blk00000001_sig00000b83 : STD_LOGIC; 
  signal blk00000001_sig00000b82 : STD_LOGIC; 
  signal blk00000001_sig00000b81 : STD_LOGIC; 
  signal blk00000001_sig00000b80 : STD_LOGIC; 
  signal blk00000001_sig00000b7f : STD_LOGIC; 
  signal blk00000001_sig00000b7e : STD_LOGIC; 
  signal blk00000001_sig00000b7d : STD_LOGIC; 
  signal blk00000001_sig00000b7c : STD_LOGIC; 
  signal blk00000001_sig00000b7b : STD_LOGIC; 
  signal blk00000001_sig00000b7a : STD_LOGIC; 
  signal blk00000001_sig00000b79 : STD_LOGIC; 
  signal blk00000001_sig00000b78 : STD_LOGIC; 
  signal blk00000001_sig00000b77 : STD_LOGIC; 
  signal blk00000001_sig00000b76 : STD_LOGIC; 
  signal blk00000001_sig00000b75 : STD_LOGIC; 
  signal blk00000001_sig00000b74 : STD_LOGIC; 
  signal blk00000001_sig00000b73 : STD_LOGIC; 
  signal blk00000001_sig00000b72 : STD_LOGIC; 
  signal blk00000001_sig00000b71 : STD_LOGIC; 
  signal blk00000001_sig00000b70 : STD_LOGIC; 
  signal blk00000001_sig00000b6f : STD_LOGIC; 
  signal blk00000001_sig00000b6e : STD_LOGIC; 
  signal blk00000001_sig00000b6d : STD_LOGIC; 
  signal blk00000001_sig00000b6c : STD_LOGIC; 
  signal blk00000001_sig00000b6b : STD_LOGIC; 
  signal blk00000001_sig00000b6a : STD_LOGIC; 
  signal blk00000001_sig00000b69 : STD_LOGIC; 
  signal blk00000001_sig00000b68 : STD_LOGIC; 
  signal blk00000001_sig00000b67 : STD_LOGIC; 
  signal blk00000001_sig00000b66 : STD_LOGIC; 
  signal blk00000001_sig00000b65 : STD_LOGIC; 
  signal blk00000001_sig00000b64 : STD_LOGIC; 
  signal blk00000001_sig00000b63 : STD_LOGIC; 
  signal blk00000001_sig00000b62 : STD_LOGIC; 
  signal blk00000001_sig00000b61 : STD_LOGIC; 
  signal blk00000001_sig00000b60 : STD_LOGIC; 
  signal blk00000001_sig00000b5f : STD_LOGIC; 
  signal blk00000001_sig00000b5e : STD_LOGIC; 
  signal blk00000001_sig00000b5d : STD_LOGIC; 
  signal blk00000001_sig00000b5c : STD_LOGIC; 
  signal blk00000001_sig00000b5b : STD_LOGIC; 
  signal blk00000001_sig00000b5a : STD_LOGIC; 
  signal blk00000001_sig00000b59 : STD_LOGIC; 
  signal blk00000001_sig00000b58 : STD_LOGIC; 
  signal blk00000001_sig00000b57 : STD_LOGIC; 
  signal blk00000001_sig00000b56 : STD_LOGIC; 
  signal blk00000001_sig00000b55 : STD_LOGIC; 
  signal blk00000001_sig00000b54 : STD_LOGIC; 
  signal blk00000001_sig00000b53 : STD_LOGIC; 
  signal blk00000001_sig00000b52 : STD_LOGIC; 
  signal blk00000001_sig00000b51 : STD_LOGIC; 
  signal blk00000001_sig00000b50 : STD_LOGIC; 
  signal blk00000001_sig00000b4f : STD_LOGIC; 
  signal blk00000001_sig00000b4e : STD_LOGIC; 
  signal blk00000001_sig00000b4d : STD_LOGIC; 
  signal blk00000001_sig00000b4c : STD_LOGIC; 
  signal blk00000001_sig00000b4b : STD_LOGIC; 
  signal blk00000001_sig00000b4a : STD_LOGIC; 
  signal blk00000001_sig00000b49 : STD_LOGIC; 
  signal blk00000001_sig00000b48 : STD_LOGIC; 
  signal blk00000001_sig00000b47 : STD_LOGIC; 
  signal blk00000001_sig00000b46 : STD_LOGIC; 
  signal blk00000001_sig00000b45 : STD_LOGIC; 
  signal blk00000001_sig00000b44 : STD_LOGIC; 
  signal blk00000001_sig00000b43 : STD_LOGIC; 
  signal blk00000001_sig00000b42 : STD_LOGIC; 
  signal blk00000001_sig00000b41 : STD_LOGIC; 
  signal blk00000001_sig00000b40 : STD_LOGIC; 
  signal blk00000001_sig00000b3f : STD_LOGIC; 
  signal blk00000001_sig00000b3e : STD_LOGIC; 
  signal blk00000001_sig00000b3d : STD_LOGIC; 
  signal blk00000001_sig00000b3c : STD_LOGIC; 
  signal blk00000001_sig00000b3b : STD_LOGIC; 
  signal blk00000001_sig00000b3a : STD_LOGIC; 
  signal blk00000001_sig00000b39 : STD_LOGIC; 
  signal blk00000001_sig00000b38 : STD_LOGIC; 
  signal blk00000001_sig00000b37 : STD_LOGIC; 
  signal blk00000001_sig00000b36 : STD_LOGIC; 
  signal blk00000001_sig00000b35 : STD_LOGIC; 
  signal blk00000001_sig00000b34 : STD_LOGIC; 
  signal blk00000001_sig00000b33 : STD_LOGIC; 
  signal blk00000001_sig00000b32 : STD_LOGIC; 
  signal blk00000001_sig00000b31 : STD_LOGIC; 
  signal blk00000001_sig00000b30 : STD_LOGIC; 
  signal blk00000001_sig00000b2f : STD_LOGIC; 
  signal blk00000001_sig00000b2e : STD_LOGIC; 
  signal blk00000001_sig00000b2d : STD_LOGIC; 
  signal blk00000001_sig00000b2c : STD_LOGIC; 
  signal blk00000001_sig00000b2b : STD_LOGIC; 
  signal blk00000001_sig00000b2a : STD_LOGIC; 
  signal blk00000001_sig00000b29 : STD_LOGIC; 
  signal blk00000001_sig00000b28 : STD_LOGIC; 
  signal blk00000001_sig00000b27 : STD_LOGIC; 
  signal blk00000001_sig00000b26 : STD_LOGIC; 
  signal blk00000001_sig00000b25 : STD_LOGIC; 
  signal blk00000001_sig00000b24 : STD_LOGIC; 
  signal blk00000001_sig00000b23 : STD_LOGIC; 
  signal blk00000001_sig00000b22 : STD_LOGIC; 
  signal blk00000001_sig00000b21 : STD_LOGIC; 
  signal blk00000001_sig00000b20 : STD_LOGIC; 
  signal blk00000001_sig00000b1f : STD_LOGIC; 
  signal blk00000001_sig00000b1e : STD_LOGIC; 
  signal blk00000001_sig00000b1d : STD_LOGIC; 
  signal blk00000001_sig00000b1c : STD_LOGIC; 
  signal blk00000001_sig00000b1b : STD_LOGIC; 
  signal blk00000001_sig00000b1a : STD_LOGIC; 
  signal blk00000001_sig00000b19 : STD_LOGIC; 
  signal blk00000001_sig00000b18 : STD_LOGIC; 
  signal blk00000001_sig00000b17 : STD_LOGIC; 
  signal blk00000001_sig00000b16 : STD_LOGIC; 
  signal blk00000001_sig00000b15 : STD_LOGIC; 
  signal blk00000001_sig00000b14 : STD_LOGIC; 
  signal blk00000001_sig00000b13 : STD_LOGIC; 
  signal blk00000001_sig00000b12 : STD_LOGIC; 
  signal blk00000001_sig00000b11 : STD_LOGIC; 
  signal blk00000001_sig00000b10 : STD_LOGIC; 
  signal blk00000001_sig00000b0f : STD_LOGIC; 
  signal blk00000001_sig00000b0e : STD_LOGIC; 
  signal blk00000001_sig00000b0d : STD_LOGIC; 
  signal blk00000001_sig00000b0c : STD_LOGIC; 
  signal blk00000001_sig00000b0b : STD_LOGIC; 
  signal blk00000001_sig00000b0a : STD_LOGIC; 
  signal blk00000001_sig00000b09 : STD_LOGIC; 
  signal blk00000001_sig00000b08 : STD_LOGIC; 
  signal blk00000001_sig00000b07 : STD_LOGIC; 
  signal blk00000001_sig00000b06 : STD_LOGIC; 
  signal blk00000001_sig00000b05 : STD_LOGIC; 
  signal blk00000001_sig00000b04 : STD_LOGIC; 
  signal blk00000001_sig00000b03 : STD_LOGIC; 
  signal blk00000001_sig00000b02 : STD_LOGIC; 
  signal blk00000001_sig00000b01 : STD_LOGIC; 
  signal blk00000001_sig00000b00 : STD_LOGIC; 
  signal blk00000001_sig00000aff : STD_LOGIC; 
  signal blk00000001_sig00000afe : STD_LOGIC; 
  signal blk00000001_sig00000afd : STD_LOGIC; 
  signal blk00000001_sig00000afc : STD_LOGIC; 
  signal blk00000001_sig00000afb : STD_LOGIC; 
  signal blk00000001_sig00000afa : STD_LOGIC; 
  signal blk00000001_sig00000af9 : STD_LOGIC; 
  signal blk00000001_sig00000af8 : STD_LOGIC; 
  signal blk00000001_sig00000af7 : STD_LOGIC; 
  signal blk00000001_sig00000af6 : STD_LOGIC; 
  signal blk00000001_sig00000af5 : STD_LOGIC; 
  signal blk00000001_sig00000af4 : STD_LOGIC; 
  signal blk00000001_sig00000af3 : STD_LOGIC; 
  signal blk00000001_sig00000af2 : STD_LOGIC; 
  signal blk00000001_sig00000af1 : STD_LOGIC; 
  signal blk00000001_sig00000af0 : STD_LOGIC; 
  signal blk00000001_sig00000aef : STD_LOGIC; 
  signal blk00000001_sig00000aee : STD_LOGIC; 
  signal blk00000001_sig00000aed : STD_LOGIC; 
  signal blk00000001_sig00000aec : STD_LOGIC; 
  signal blk00000001_sig00000aeb : STD_LOGIC; 
  signal blk00000001_sig00000aea : STD_LOGIC; 
  signal blk00000001_sig00000ae9 : STD_LOGIC; 
  signal blk00000001_sig00000ae8 : STD_LOGIC; 
  signal blk00000001_sig00000ae7 : STD_LOGIC; 
  signal blk00000001_sig00000ae6 : STD_LOGIC; 
  signal blk00000001_sig00000ae5 : STD_LOGIC; 
  signal blk00000001_sig00000ae4 : STD_LOGIC; 
  signal blk00000001_sig00000ae3 : STD_LOGIC; 
  signal blk00000001_sig00000ae2 : STD_LOGIC; 
  signal blk00000001_sig00000ae1 : STD_LOGIC; 
  signal blk00000001_sig00000ae0 : STD_LOGIC; 
  signal blk00000001_sig00000adf : STD_LOGIC; 
  signal blk00000001_sig00000ade : STD_LOGIC; 
  signal blk00000001_sig00000add : STD_LOGIC; 
  signal blk00000001_sig00000adc : STD_LOGIC; 
  signal blk00000001_sig00000adb : STD_LOGIC; 
  signal blk00000001_sig00000ada : STD_LOGIC; 
  signal blk00000001_sig00000ad9 : STD_LOGIC; 
  signal blk00000001_sig00000ad8 : STD_LOGIC; 
  signal blk00000001_sig00000ad7 : STD_LOGIC; 
  signal blk00000001_sig00000ad6 : STD_LOGIC; 
  signal blk00000001_sig00000ad5 : STD_LOGIC; 
  signal blk00000001_sig00000ad4 : STD_LOGIC; 
  signal blk00000001_sig00000ad3 : STD_LOGIC; 
  signal blk00000001_sig00000ad2 : STD_LOGIC; 
  signal blk00000001_sig00000ad1 : STD_LOGIC; 
  signal blk00000001_sig00000ad0 : STD_LOGIC; 
  signal blk00000001_sig00000acf : STD_LOGIC; 
  signal blk00000001_sig00000ace : STD_LOGIC; 
  signal blk00000001_sig00000acd : STD_LOGIC; 
  signal blk00000001_sig00000acc : STD_LOGIC; 
  signal blk00000001_sig00000acb : STD_LOGIC; 
  signal blk00000001_sig00000aca : STD_LOGIC; 
  signal blk00000001_sig00000ac9 : STD_LOGIC; 
  signal blk00000001_sig00000ac8 : STD_LOGIC; 
  signal blk00000001_sig00000ac7 : STD_LOGIC; 
  signal blk00000001_sig00000ac6 : STD_LOGIC; 
  signal blk00000001_sig00000ac5 : STD_LOGIC; 
  signal blk00000001_sig00000ac4 : STD_LOGIC; 
  signal blk00000001_sig00000ac3 : STD_LOGIC; 
  signal blk00000001_sig00000ac2 : STD_LOGIC; 
  signal blk00000001_sig00000ac1 : STD_LOGIC; 
  signal blk00000001_sig00000ac0 : STD_LOGIC; 
  signal blk00000001_sig00000abf : STD_LOGIC; 
  signal blk00000001_sig00000abe : STD_LOGIC; 
  signal blk00000001_sig00000abd : STD_LOGIC; 
  signal blk00000001_sig00000abc : STD_LOGIC; 
  signal blk00000001_sig00000abb : STD_LOGIC; 
  signal blk00000001_sig00000aba : STD_LOGIC; 
  signal blk00000001_sig00000ab9 : STD_LOGIC; 
  signal blk00000001_sig00000ab8 : STD_LOGIC; 
  signal blk00000001_sig00000ab7 : STD_LOGIC; 
  signal blk00000001_sig00000ab6 : STD_LOGIC; 
  signal blk00000001_sig00000ab5 : STD_LOGIC; 
  signal blk00000001_sig00000ab4 : STD_LOGIC; 
  signal blk00000001_sig00000ab3 : STD_LOGIC; 
  signal blk00000001_sig00000ab2 : STD_LOGIC; 
  signal blk00000001_sig00000ab1 : STD_LOGIC; 
  signal blk00000001_sig00000ab0 : STD_LOGIC; 
  signal blk00000001_sig00000aaf : STD_LOGIC; 
  signal blk00000001_sig00000aae : STD_LOGIC; 
  signal blk00000001_sig00000aad : STD_LOGIC; 
  signal blk00000001_sig00000aac : STD_LOGIC; 
  signal blk00000001_sig00000aab : STD_LOGIC; 
  signal blk00000001_sig00000aaa : STD_LOGIC; 
  signal blk00000001_sig00000aa9 : STD_LOGIC; 
  signal blk00000001_sig00000aa8 : STD_LOGIC; 
  signal blk00000001_sig00000aa7 : STD_LOGIC; 
  signal blk00000001_sig00000aa6 : STD_LOGIC; 
  signal blk00000001_sig00000aa5 : STD_LOGIC; 
  signal blk00000001_sig00000aa4 : STD_LOGIC; 
  signal blk00000001_sig00000aa3 : STD_LOGIC; 
  signal blk00000001_sig00000aa2 : STD_LOGIC; 
  signal blk00000001_sig00000aa1 : STD_LOGIC; 
  signal blk00000001_sig00000aa0 : STD_LOGIC; 
  signal blk00000001_sig00000a9f : STD_LOGIC; 
  signal blk00000001_sig00000a9e : STD_LOGIC; 
  signal blk00000001_sig00000a9d : STD_LOGIC; 
  signal blk00000001_sig00000a9c : STD_LOGIC; 
  signal blk00000001_sig00000a9b : STD_LOGIC; 
  signal blk00000001_sig00000a9a : STD_LOGIC; 
  signal blk00000001_sig00000a99 : STD_LOGIC; 
  signal blk00000001_sig00000a98 : STD_LOGIC; 
  signal blk00000001_sig00000a97 : STD_LOGIC; 
  signal blk00000001_sig00000a96 : STD_LOGIC; 
  signal blk00000001_sig00000a95 : STD_LOGIC; 
  signal blk00000001_sig00000a94 : STD_LOGIC; 
  signal blk00000001_sig00000a93 : STD_LOGIC; 
  signal blk00000001_sig00000a92 : STD_LOGIC; 
  signal blk00000001_sig00000a91 : STD_LOGIC; 
  signal blk00000001_sig00000a90 : STD_LOGIC; 
  signal blk00000001_sig00000a8f : STD_LOGIC; 
  signal blk00000001_sig00000a8e : STD_LOGIC; 
  signal blk00000001_sig00000a8d : STD_LOGIC; 
  signal blk00000001_sig00000a8c : STD_LOGIC; 
  signal blk00000001_sig00000a8b : STD_LOGIC; 
  signal blk00000001_sig00000a8a : STD_LOGIC; 
  signal blk00000001_sig00000a89 : STD_LOGIC; 
  signal blk00000001_sig00000a88 : STD_LOGIC; 
  signal blk00000001_sig00000a87 : STD_LOGIC; 
  signal blk00000001_sig00000a86 : STD_LOGIC; 
  signal blk00000001_sig00000a85 : STD_LOGIC; 
  signal blk00000001_sig00000a84 : STD_LOGIC; 
  signal blk00000001_sig00000a83 : STD_LOGIC; 
  signal blk00000001_sig00000a82 : STD_LOGIC; 
  signal blk00000001_sig00000a81 : STD_LOGIC; 
  signal blk00000001_sig00000a80 : STD_LOGIC; 
  signal blk00000001_sig00000a7f : STD_LOGIC; 
  signal blk00000001_sig00000a7e : STD_LOGIC; 
  signal blk00000001_sig00000a7d : STD_LOGIC; 
  signal blk00000001_sig00000a7c : STD_LOGIC; 
  signal blk00000001_sig00000a7b : STD_LOGIC; 
  signal blk00000001_sig00000a7a : STD_LOGIC; 
  signal blk00000001_sig00000a79 : STD_LOGIC; 
  signal blk00000001_sig00000a78 : STD_LOGIC; 
  signal blk00000001_sig00000a77 : STD_LOGIC; 
  signal blk00000001_sig00000a76 : STD_LOGIC; 
  signal blk00000001_sig00000a75 : STD_LOGIC; 
  signal blk00000001_sig00000a74 : STD_LOGIC; 
  signal blk00000001_sig00000a73 : STD_LOGIC; 
  signal blk00000001_sig00000a72 : STD_LOGIC; 
  signal blk00000001_sig00000a71 : STD_LOGIC; 
  signal blk00000001_sig00000a70 : STD_LOGIC; 
  signal blk00000001_sig00000a6f : STD_LOGIC; 
  signal blk00000001_sig00000a6e : STD_LOGIC; 
  signal blk00000001_sig00000a6d : STD_LOGIC; 
  signal blk00000001_sig00000a6c : STD_LOGIC; 
  signal blk00000001_sig00000a6b : STD_LOGIC; 
  signal blk00000001_sig00000a6a : STD_LOGIC; 
  signal blk00000001_sig00000a69 : STD_LOGIC; 
  signal blk00000001_sig00000a68 : STD_LOGIC; 
  signal blk00000001_sig00000a67 : STD_LOGIC; 
  signal blk00000001_sig00000a66 : STD_LOGIC; 
  signal blk00000001_sig00000a65 : STD_LOGIC; 
  signal blk00000001_sig00000a64 : STD_LOGIC; 
  signal blk00000001_sig00000a63 : STD_LOGIC; 
  signal blk00000001_sig00000a62 : STD_LOGIC; 
  signal blk00000001_sig00000a61 : STD_LOGIC; 
  signal blk00000001_sig00000a60 : STD_LOGIC; 
  signal blk00000001_sig00000a5f : STD_LOGIC; 
  signal blk00000001_sig00000a5e : STD_LOGIC; 
  signal blk00000001_sig00000a5d : STD_LOGIC; 
  signal blk00000001_sig00000a5c : STD_LOGIC; 
  signal blk00000001_sig00000a5b : STD_LOGIC; 
  signal blk00000001_sig00000a5a : STD_LOGIC; 
  signal blk00000001_sig00000a59 : STD_LOGIC; 
  signal blk00000001_sig00000a58 : STD_LOGIC; 
  signal blk00000001_sig00000a57 : STD_LOGIC; 
  signal blk00000001_sig00000a56 : STD_LOGIC; 
  signal blk00000001_sig00000a55 : STD_LOGIC; 
  signal blk00000001_sig00000a54 : STD_LOGIC; 
  signal blk00000001_sig00000a53 : STD_LOGIC; 
  signal blk00000001_sig00000a52 : STD_LOGIC; 
  signal blk00000001_sig00000a51 : STD_LOGIC; 
  signal blk00000001_sig00000a50 : STD_LOGIC; 
  signal blk00000001_sig00000a4f : STD_LOGIC; 
  signal blk00000001_sig00000a4e : STD_LOGIC; 
  signal blk00000001_sig00000a4d : STD_LOGIC; 
  signal blk00000001_sig00000a4c : STD_LOGIC; 
  signal blk00000001_sig00000a4b : STD_LOGIC; 
  signal blk00000001_sig00000a4a : STD_LOGIC; 
  signal blk00000001_sig00000a49 : STD_LOGIC; 
  signal blk00000001_sig00000a48 : STD_LOGIC; 
  signal blk00000001_sig00000a47 : STD_LOGIC; 
  signal blk00000001_sig00000a46 : STD_LOGIC; 
  signal blk00000001_sig00000a45 : STD_LOGIC; 
  signal blk00000001_sig00000a44 : STD_LOGIC; 
  signal blk00000001_sig00000a43 : STD_LOGIC; 
  signal blk00000001_sig00000a42 : STD_LOGIC; 
  signal blk00000001_sig00000a41 : STD_LOGIC; 
  signal blk00000001_sig00000a40 : STD_LOGIC; 
  signal blk00000001_sig00000a3f : STD_LOGIC; 
  signal blk00000001_sig00000a3e : STD_LOGIC; 
  signal blk00000001_sig00000a3d : STD_LOGIC; 
  signal blk00000001_sig00000a3c : STD_LOGIC; 
  signal blk00000001_sig00000a3b : STD_LOGIC; 
  signal blk00000001_sig00000a3a : STD_LOGIC; 
  signal blk00000001_sig00000a39 : STD_LOGIC; 
  signal blk00000001_sig00000a38 : STD_LOGIC; 
  signal blk00000001_sig00000a37 : STD_LOGIC; 
  signal blk00000001_sig00000a36 : STD_LOGIC; 
  signal blk00000001_sig00000a35 : STD_LOGIC; 
  signal blk00000001_sig00000a34 : STD_LOGIC; 
  signal blk00000001_sig00000a33 : STD_LOGIC; 
  signal blk00000001_sig00000a32 : STD_LOGIC; 
  signal blk00000001_sig00000a31 : STD_LOGIC; 
  signal blk00000001_sig00000a30 : STD_LOGIC; 
  signal blk00000001_sig00000a2f : STD_LOGIC; 
  signal blk00000001_sig00000a2e : STD_LOGIC; 
  signal blk00000001_sig00000a2d : STD_LOGIC; 
  signal blk00000001_sig00000a2c : STD_LOGIC; 
  signal blk00000001_sig00000a2b : STD_LOGIC; 
  signal blk00000001_sig00000a2a : STD_LOGIC; 
  signal blk00000001_sig00000a29 : STD_LOGIC; 
  signal blk00000001_sig00000a28 : STD_LOGIC; 
  signal blk00000001_sig00000a27 : STD_LOGIC; 
  signal blk00000001_sig00000a26 : STD_LOGIC; 
  signal blk00000001_sig00000a25 : STD_LOGIC; 
  signal blk00000001_sig00000a24 : STD_LOGIC; 
  signal blk00000001_sig00000a23 : STD_LOGIC; 
  signal blk00000001_sig00000a22 : STD_LOGIC; 
  signal blk00000001_sig00000a21 : STD_LOGIC; 
  signal blk00000001_sig00000a20 : STD_LOGIC; 
  signal blk00000001_sig00000a1f : STD_LOGIC; 
  signal blk00000001_sig00000a1e : STD_LOGIC; 
  signal blk00000001_sig00000a1d : STD_LOGIC; 
  signal blk00000001_sig00000a1c : STD_LOGIC; 
  signal blk00000001_sig00000a1b : STD_LOGIC; 
  signal blk00000001_sig00000a1a : STD_LOGIC; 
  signal blk00000001_sig00000a19 : STD_LOGIC; 
  signal blk00000001_sig00000a18 : STD_LOGIC; 
  signal blk00000001_sig00000a17 : STD_LOGIC; 
  signal blk00000001_sig00000a16 : STD_LOGIC; 
  signal blk00000001_sig00000a15 : STD_LOGIC; 
  signal blk00000001_sig00000a14 : STD_LOGIC; 
  signal blk00000001_sig00000a13 : STD_LOGIC; 
  signal blk00000001_sig00000a12 : STD_LOGIC; 
  signal blk00000001_sig00000a11 : STD_LOGIC; 
  signal blk00000001_sig00000a10 : STD_LOGIC; 
  signal blk00000001_sig00000a0f : STD_LOGIC; 
  signal blk00000001_sig00000a0e : STD_LOGIC; 
  signal blk00000001_sig00000a0d : STD_LOGIC; 
  signal blk00000001_sig00000a0c : STD_LOGIC; 
  signal blk00000001_sig00000a0b : STD_LOGIC; 
  signal blk00000001_sig00000a0a : STD_LOGIC; 
  signal blk00000001_sig00000a09 : STD_LOGIC; 
  signal blk00000001_sig00000a08 : STD_LOGIC; 
  signal blk00000001_sig00000a07 : STD_LOGIC; 
  signal blk00000001_sig00000a06 : STD_LOGIC; 
  signal blk00000001_sig00000a05 : STD_LOGIC; 
  signal blk00000001_sig00000a04 : STD_LOGIC; 
  signal blk00000001_sig00000a03 : STD_LOGIC; 
  signal blk00000001_sig00000a02 : STD_LOGIC; 
  signal blk00000001_sig00000a01 : STD_LOGIC; 
  signal blk00000001_sig00000a00 : STD_LOGIC; 
  signal blk00000001_sig000009ff : STD_LOGIC; 
  signal blk00000001_sig000009fe : STD_LOGIC; 
  signal blk00000001_sig000009fd : STD_LOGIC; 
  signal blk00000001_sig000009fc : STD_LOGIC; 
  signal blk00000001_sig000009fb : STD_LOGIC; 
  signal blk00000001_sig000009fa : STD_LOGIC; 
  signal blk00000001_sig000009f9 : STD_LOGIC; 
  signal blk00000001_sig000009f8 : STD_LOGIC; 
  signal blk00000001_sig000009f7 : STD_LOGIC; 
  signal blk00000001_sig000009f6 : STD_LOGIC; 
  signal blk00000001_sig000009f5 : STD_LOGIC; 
  signal blk00000001_sig000009f4 : STD_LOGIC; 
  signal blk00000001_sig000009f3 : STD_LOGIC; 
  signal blk00000001_sig000009f2 : STD_LOGIC; 
  signal blk00000001_sig000009f1 : STD_LOGIC; 
  signal blk00000001_sig000009f0 : STD_LOGIC; 
  signal blk00000001_sig000009ef : STD_LOGIC; 
  signal blk00000001_sig000009ee : STD_LOGIC; 
  signal blk00000001_sig000009ed : STD_LOGIC; 
  signal blk00000001_sig000009ec : STD_LOGIC; 
  signal blk00000001_sig000009eb : STD_LOGIC; 
  signal blk00000001_sig000009ea : STD_LOGIC; 
  signal blk00000001_sig000009e9 : STD_LOGIC; 
  signal blk00000001_sig000009e8 : STD_LOGIC; 
  signal blk00000001_sig000009e7 : STD_LOGIC; 
  signal blk00000001_sig000009e6 : STD_LOGIC; 
  signal blk00000001_sig000009e5 : STD_LOGIC; 
  signal blk00000001_sig000009e4 : STD_LOGIC; 
  signal blk00000001_sig000009e3 : STD_LOGIC; 
  signal blk00000001_sig000009e2 : STD_LOGIC; 
  signal blk00000001_sig000009e1 : STD_LOGIC; 
  signal blk00000001_sig000009e0 : STD_LOGIC; 
  signal blk00000001_sig000009df : STD_LOGIC; 
  signal blk00000001_sig000009de : STD_LOGIC; 
  signal blk00000001_sig000009dd : STD_LOGIC; 
  signal blk00000001_sig000009dc : STD_LOGIC; 
  signal blk00000001_sig000009db : STD_LOGIC; 
  signal blk00000001_sig000009da : STD_LOGIC; 
  signal blk00000001_sig000009d9 : STD_LOGIC; 
  signal blk00000001_sig000009d8 : STD_LOGIC; 
  signal blk00000001_sig000009d7 : STD_LOGIC; 
  signal blk00000001_sig000009d6 : STD_LOGIC; 
  signal blk00000001_sig000009d5 : STD_LOGIC; 
  signal blk00000001_sig000009d4 : STD_LOGIC; 
  signal blk00000001_sig000009d3 : STD_LOGIC; 
  signal blk00000001_sig000009d2 : STD_LOGIC; 
  signal blk00000001_sig000009d1 : STD_LOGIC; 
  signal blk00000001_sig000009d0 : STD_LOGIC; 
  signal blk00000001_sig000009cf : STD_LOGIC; 
  signal blk00000001_sig000009ce : STD_LOGIC; 
  signal blk00000001_sig000009cd : STD_LOGIC; 
  signal blk00000001_sig000009cc : STD_LOGIC; 
  signal blk00000001_sig000009cb : STD_LOGIC; 
  signal blk00000001_sig000009ca : STD_LOGIC; 
  signal blk00000001_sig000009c9 : STD_LOGIC; 
  signal blk00000001_sig000009c8 : STD_LOGIC; 
  signal blk00000001_sig000009c7 : STD_LOGIC; 
  signal blk00000001_sig000009c6 : STD_LOGIC; 
  signal blk00000001_sig000009c5 : STD_LOGIC; 
  signal blk00000001_sig000009c4 : STD_LOGIC; 
  signal blk00000001_sig000009c3 : STD_LOGIC; 
  signal blk00000001_sig000009c2 : STD_LOGIC; 
  signal blk00000001_sig000009c1 : STD_LOGIC; 
  signal blk00000001_sig000009c0 : STD_LOGIC; 
  signal blk00000001_sig000009bf : STD_LOGIC; 
  signal blk00000001_sig000009be : STD_LOGIC; 
  signal blk00000001_sig000009bd : STD_LOGIC; 
  signal blk00000001_sig000009bc : STD_LOGIC; 
  signal blk00000001_sig000009bb : STD_LOGIC; 
  signal blk00000001_sig000009ba : STD_LOGIC; 
  signal blk00000001_sig000009b9 : STD_LOGIC; 
  signal blk00000001_sig000009b8 : STD_LOGIC; 
  signal blk00000001_sig000009b7 : STD_LOGIC; 
  signal blk00000001_sig000009b6 : STD_LOGIC; 
  signal blk00000001_sig000009b5 : STD_LOGIC; 
  signal blk00000001_sig000009b4 : STD_LOGIC; 
  signal blk00000001_sig000009b3 : STD_LOGIC; 
  signal blk00000001_sig000009b2 : STD_LOGIC; 
  signal blk00000001_sig000009b1 : STD_LOGIC; 
  signal blk00000001_sig000009b0 : STD_LOGIC; 
  signal blk00000001_sig000009af : STD_LOGIC; 
  signal blk00000001_sig000009ae : STD_LOGIC; 
  signal blk00000001_sig000009ad : STD_LOGIC; 
  signal blk00000001_sig000009ac : STD_LOGIC; 
  signal blk00000001_sig000009ab : STD_LOGIC; 
  signal blk00000001_sig000009aa : STD_LOGIC; 
  signal blk00000001_sig000009a9 : STD_LOGIC; 
  signal blk00000001_sig000009a8 : STD_LOGIC; 
  signal blk00000001_sig000009a7 : STD_LOGIC; 
  signal blk00000001_sig000009a6 : STD_LOGIC; 
  signal blk00000001_sig000009a5 : STD_LOGIC; 
  signal blk00000001_sig000009a4 : STD_LOGIC; 
  signal blk00000001_sig000009a3 : STD_LOGIC; 
  signal blk00000001_sig000009a2 : STD_LOGIC; 
  signal blk00000001_sig000009a1 : STD_LOGIC; 
  signal blk00000001_sig000009a0 : STD_LOGIC; 
  signal blk00000001_sig0000099f : STD_LOGIC; 
  signal blk00000001_sig0000099e : STD_LOGIC; 
  signal blk00000001_sig0000099d : STD_LOGIC; 
  signal blk00000001_sig0000099c : STD_LOGIC; 
  signal blk00000001_sig0000099b : STD_LOGIC; 
  signal blk00000001_sig0000099a : STD_LOGIC; 
  signal blk00000001_sig00000999 : STD_LOGIC; 
  signal blk00000001_sig00000998 : STD_LOGIC; 
  signal blk00000001_sig00000997 : STD_LOGIC; 
  signal blk00000001_sig00000996 : STD_LOGIC; 
  signal blk00000001_sig00000995 : STD_LOGIC; 
  signal blk00000001_sig00000994 : STD_LOGIC; 
  signal blk00000001_sig00000993 : STD_LOGIC; 
  signal blk00000001_sig00000992 : STD_LOGIC; 
  signal blk00000001_sig00000991 : STD_LOGIC; 
  signal blk00000001_sig00000990 : STD_LOGIC; 
  signal blk00000001_sig0000098f : STD_LOGIC; 
  signal blk00000001_sig0000098e : STD_LOGIC; 
  signal blk00000001_sig0000098d : STD_LOGIC; 
  signal blk00000001_sig0000098c : STD_LOGIC; 
  signal blk00000001_sig0000098b : STD_LOGIC; 
  signal blk00000001_sig0000098a : STD_LOGIC; 
  signal blk00000001_sig00000989 : STD_LOGIC; 
  signal blk00000001_sig00000988 : STD_LOGIC; 
  signal blk00000001_sig00000987 : STD_LOGIC; 
  signal blk00000001_sig00000986 : STD_LOGIC; 
  signal blk00000001_sig00000985 : STD_LOGIC; 
  signal blk00000001_sig00000984 : STD_LOGIC; 
  signal blk00000001_sig00000983 : STD_LOGIC; 
  signal blk00000001_sig00000982 : STD_LOGIC; 
  signal blk00000001_sig00000981 : STD_LOGIC; 
  signal blk00000001_sig00000980 : STD_LOGIC; 
  signal blk00000001_sig0000097f : STD_LOGIC; 
  signal blk00000001_sig0000097e : STD_LOGIC; 
  signal blk00000001_sig0000097d : STD_LOGIC; 
  signal blk00000001_sig0000097c : STD_LOGIC; 
  signal blk00000001_sig0000097b : STD_LOGIC; 
  signal blk00000001_sig0000097a : STD_LOGIC; 
  signal blk00000001_sig00000979 : STD_LOGIC; 
  signal blk00000001_sig00000978 : STD_LOGIC; 
  signal blk00000001_sig00000977 : STD_LOGIC; 
  signal blk00000001_sig00000976 : STD_LOGIC; 
  signal blk00000001_sig00000975 : STD_LOGIC; 
  signal blk00000001_sig00000974 : STD_LOGIC; 
  signal blk00000001_sig00000973 : STD_LOGIC; 
  signal blk00000001_sig00000972 : STD_LOGIC; 
  signal blk00000001_sig00000971 : STD_LOGIC; 
  signal blk00000001_sig00000970 : STD_LOGIC; 
  signal blk00000001_sig0000096f : STD_LOGIC; 
  signal blk00000001_sig0000096e : STD_LOGIC; 
  signal blk00000001_sig0000096d : STD_LOGIC; 
  signal blk00000001_sig0000096c : STD_LOGIC; 
  signal blk00000001_sig0000096b : STD_LOGIC; 
  signal blk00000001_sig0000096a : STD_LOGIC; 
  signal blk00000001_sig00000969 : STD_LOGIC; 
  signal blk00000001_sig00000968 : STD_LOGIC; 
  signal blk00000001_sig00000967 : STD_LOGIC; 
  signal blk00000001_sig00000966 : STD_LOGIC; 
  signal blk00000001_sig00000965 : STD_LOGIC; 
  signal blk00000001_sig00000964 : STD_LOGIC; 
  signal blk00000001_sig00000963 : STD_LOGIC; 
  signal blk00000001_sig00000962 : STD_LOGIC; 
  signal blk00000001_sig00000961 : STD_LOGIC; 
  signal blk00000001_sig00000960 : STD_LOGIC; 
  signal blk00000001_sig0000095f : STD_LOGIC; 
  signal blk00000001_sig0000095e : STD_LOGIC; 
  signal blk00000001_sig0000095d : STD_LOGIC; 
  signal blk00000001_sig0000095c : STD_LOGIC; 
  signal blk00000001_sig0000095b : STD_LOGIC; 
  signal blk00000001_sig0000095a : STD_LOGIC; 
  signal blk00000001_sig00000959 : STD_LOGIC; 
  signal blk00000001_sig00000958 : STD_LOGIC; 
  signal blk00000001_sig00000957 : STD_LOGIC; 
  signal blk00000001_sig00000956 : STD_LOGIC; 
  signal blk00000001_sig00000955 : STD_LOGIC; 
  signal blk00000001_sig00000954 : STD_LOGIC; 
  signal blk00000001_sig00000953 : STD_LOGIC; 
  signal blk00000001_sig00000952 : STD_LOGIC; 
  signal blk00000001_sig00000951 : STD_LOGIC; 
  signal blk00000001_sig00000950 : STD_LOGIC; 
  signal blk00000001_sig0000094f : STD_LOGIC; 
  signal blk00000001_sig0000094e : STD_LOGIC; 
  signal blk00000001_sig0000094d : STD_LOGIC; 
  signal blk00000001_sig0000094c : STD_LOGIC; 
  signal blk00000001_sig0000094b : STD_LOGIC; 
  signal blk00000001_sig0000094a : STD_LOGIC; 
  signal blk00000001_sig00000949 : STD_LOGIC; 
  signal blk00000001_sig00000948 : STD_LOGIC; 
  signal blk00000001_sig00000947 : STD_LOGIC; 
  signal blk00000001_sig00000946 : STD_LOGIC; 
  signal blk00000001_sig00000945 : STD_LOGIC; 
  signal blk00000001_sig00000944 : STD_LOGIC; 
  signal blk00000001_sig00000943 : STD_LOGIC; 
  signal blk00000001_sig00000942 : STD_LOGIC; 
  signal blk00000001_sig00000941 : STD_LOGIC; 
  signal blk00000001_sig00000940 : STD_LOGIC; 
  signal blk00000001_sig0000093f : STD_LOGIC; 
  signal blk00000001_sig0000093e : STD_LOGIC; 
  signal blk00000001_sig0000093d : STD_LOGIC; 
  signal blk00000001_sig0000093c : STD_LOGIC; 
  signal blk00000001_sig0000093b : STD_LOGIC; 
  signal blk00000001_sig0000093a : STD_LOGIC; 
  signal blk00000001_sig00000939 : STD_LOGIC; 
  signal blk00000001_sig00000938 : STD_LOGIC; 
  signal blk00000001_sig00000937 : STD_LOGIC; 
  signal blk00000001_sig00000936 : STD_LOGIC; 
  signal blk00000001_sig00000935 : STD_LOGIC; 
  signal blk00000001_sig00000934 : STD_LOGIC; 
  signal blk00000001_sig00000933 : STD_LOGIC; 
  signal blk00000001_sig00000932 : STD_LOGIC; 
  signal blk00000001_sig00000931 : STD_LOGIC; 
  signal blk00000001_sig00000930 : STD_LOGIC; 
  signal blk00000001_sig0000092f : STD_LOGIC; 
  signal blk00000001_sig0000092e : STD_LOGIC; 
  signal blk00000001_sig0000092d : STD_LOGIC; 
  signal blk00000001_sig0000092c : STD_LOGIC; 
  signal blk00000001_sig0000092b : STD_LOGIC; 
  signal blk00000001_sig0000092a : STD_LOGIC; 
  signal blk00000001_sig00000929 : STD_LOGIC; 
  signal blk00000001_sig00000928 : STD_LOGIC; 
  signal blk00000001_sig00000927 : STD_LOGIC; 
  signal blk00000001_sig00000926 : STD_LOGIC; 
  signal blk00000001_sig00000925 : STD_LOGIC; 
  signal blk00000001_sig00000924 : STD_LOGIC; 
  signal blk00000001_sig00000922 : STD_LOGIC; 
  signal blk00000001_sig00000921 : STD_LOGIC; 
  signal blk00000001_sig00000920 : STD_LOGIC; 
  signal blk00000001_sig0000091f : STD_LOGIC; 
  signal blk00000001_sig0000091e : STD_LOGIC; 
  signal blk00000001_sig0000091d : STD_LOGIC; 
  signal blk00000001_sig0000091c : STD_LOGIC; 
  signal blk00000001_sig0000091b : STD_LOGIC; 
  signal blk00000001_sig0000091a : STD_LOGIC; 
  signal blk00000001_sig00000919 : STD_LOGIC; 
  signal blk00000001_sig00000918 : STD_LOGIC; 
  signal blk00000001_sig00000917 : STD_LOGIC; 
  signal blk00000001_sig00000916 : STD_LOGIC; 
  signal blk00000001_sig00000915 : STD_LOGIC; 
  signal blk00000001_sig00000914 : STD_LOGIC; 
  signal blk00000001_sig00000913 : STD_LOGIC; 
  signal blk00000001_sig00000912 : STD_LOGIC; 
  signal blk00000001_sig00000911 : STD_LOGIC; 
  signal blk00000001_sig00000910 : STD_LOGIC; 
  signal blk00000001_sig0000090f : STD_LOGIC; 
  signal blk00000001_sig0000090e : STD_LOGIC; 
  signal blk00000001_sig0000090d : STD_LOGIC; 
  signal blk00000001_sig0000090c : STD_LOGIC; 
  signal blk00000001_sig0000090b : STD_LOGIC; 
  signal blk00000001_sig0000090a : STD_LOGIC; 
  signal blk00000001_sig00000909 : STD_LOGIC; 
  signal blk00000001_sig00000908 : STD_LOGIC; 
  signal blk00000001_sig00000907 : STD_LOGIC; 
  signal blk00000001_sig00000906 : STD_LOGIC; 
  signal blk00000001_sig00000905 : STD_LOGIC; 
  signal blk00000001_sig00000904 : STD_LOGIC; 
  signal blk00000001_sig00000903 : STD_LOGIC; 
  signal blk00000001_sig00000902 : STD_LOGIC; 
  signal blk00000001_sig00000901 : STD_LOGIC; 
  signal blk00000001_sig00000900 : STD_LOGIC; 
  signal blk00000001_sig000008ff : STD_LOGIC; 
  signal blk00000001_sig000008fe : STD_LOGIC; 
  signal blk00000001_sig000008fd : STD_LOGIC; 
  signal blk00000001_sig000008fc : STD_LOGIC; 
  signal blk00000001_sig000008fb : STD_LOGIC; 
  signal blk00000001_sig000008fa : STD_LOGIC; 
  signal blk00000001_sig000008f9 : STD_LOGIC; 
  signal blk00000001_sig000008f8 : STD_LOGIC; 
  signal blk00000001_sig000008f7 : STD_LOGIC; 
  signal blk00000001_sig000008f6 : STD_LOGIC; 
  signal blk00000001_sig000008f5 : STD_LOGIC; 
  signal blk00000001_sig000008f4 : STD_LOGIC; 
  signal blk00000001_sig000008f3 : STD_LOGIC; 
  signal blk00000001_sig000008f2 : STD_LOGIC; 
  signal blk00000001_sig000008f1 : STD_LOGIC; 
  signal blk00000001_sig000008f0 : STD_LOGIC; 
  signal blk00000001_sig000008ef : STD_LOGIC; 
  signal blk00000001_sig000008ee : STD_LOGIC; 
  signal blk00000001_sig000008ed : STD_LOGIC; 
  signal blk00000001_sig000008ec : STD_LOGIC; 
  signal blk00000001_sig000008eb : STD_LOGIC; 
  signal blk00000001_sig000008ea : STD_LOGIC; 
  signal blk00000001_sig000008e9 : STD_LOGIC; 
  signal blk00000001_sig000008e8 : STD_LOGIC; 
  signal blk00000001_sig000008e7 : STD_LOGIC; 
  signal blk00000001_sig000008e6 : STD_LOGIC; 
  signal blk00000001_sig000008e5 : STD_LOGIC; 
  signal blk00000001_sig000008e4 : STD_LOGIC; 
  signal blk00000001_sig000008e3 : STD_LOGIC; 
  signal blk00000001_sig000008e2 : STD_LOGIC; 
  signal blk00000001_sig000008e1 : STD_LOGIC; 
  signal blk00000001_sig000008e0 : STD_LOGIC; 
  signal blk00000001_sig000008df : STD_LOGIC; 
  signal blk00000001_sig000008de : STD_LOGIC; 
  signal blk00000001_sig000008dd : STD_LOGIC; 
  signal blk00000001_sig000008dc : STD_LOGIC; 
  signal blk00000001_sig000008db : STD_LOGIC; 
  signal blk00000001_sig000008da : STD_LOGIC; 
  signal blk00000001_sig000008d9 : STD_LOGIC; 
  signal blk00000001_sig000008d8 : STD_LOGIC; 
  signal blk00000001_sig000008d7 : STD_LOGIC; 
  signal blk00000001_sig000008d6 : STD_LOGIC; 
  signal blk00000001_sig000008d5 : STD_LOGIC; 
  signal blk00000001_sig000008d4 : STD_LOGIC; 
  signal blk00000001_sig000008d3 : STD_LOGIC; 
  signal blk00000001_sig000008d2 : STD_LOGIC; 
  signal blk00000001_sig000008d1 : STD_LOGIC; 
  signal blk00000001_sig000008d0 : STD_LOGIC; 
  signal blk00000001_sig000008cf : STD_LOGIC; 
  signal blk00000001_sig000008ce : STD_LOGIC; 
  signal blk00000001_sig000008cd : STD_LOGIC; 
  signal blk00000001_sig000008cc : STD_LOGIC; 
  signal blk00000001_sig000008cb : STD_LOGIC; 
  signal blk00000001_sig000008ca : STD_LOGIC; 
  signal blk00000001_sig000008c9 : STD_LOGIC; 
  signal blk00000001_sig000008c8 : STD_LOGIC; 
  signal blk00000001_sig000008c7 : STD_LOGIC; 
  signal blk00000001_sig000008c6 : STD_LOGIC; 
  signal blk00000001_sig000008c5 : STD_LOGIC; 
  signal blk00000001_sig000008c4 : STD_LOGIC; 
  signal blk00000001_sig000008c3 : STD_LOGIC; 
  signal blk00000001_sig000008c2 : STD_LOGIC; 
  signal blk00000001_sig000008c1 : STD_LOGIC; 
  signal blk00000001_sig000008c0 : STD_LOGIC; 
  signal blk00000001_sig000008bf : STD_LOGIC; 
  signal blk00000001_sig000008be : STD_LOGIC; 
  signal blk00000001_sig000008bd : STD_LOGIC; 
  signal blk00000001_sig000008bc : STD_LOGIC; 
  signal blk00000001_sig000008bb : STD_LOGIC; 
  signal blk00000001_sig000008ba : STD_LOGIC; 
  signal blk00000001_sig000008b9 : STD_LOGIC; 
  signal blk00000001_sig000008b8 : STD_LOGIC; 
  signal blk00000001_sig000008b7 : STD_LOGIC; 
  signal blk00000001_sig000008b6 : STD_LOGIC; 
  signal blk00000001_sig000008b5 : STD_LOGIC; 
  signal blk00000001_sig000008b4 : STD_LOGIC; 
  signal blk00000001_sig000008b3 : STD_LOGIC; 
  signal blk00000001_sig000008b2 : STD_LOGIC; 
  signal blk00000001_sig000008b1 : STD_LOGIC; 
  signal blk00000001_sig000008b0 : STD_LOGIC; 
  signal blk00000001_sig000008af : STD_LOGIC; 
  signal blk00000001_sig000008ae : STD_LOGIC; 
  signal blk00000001_sig000008ad : STD_LOGIC; 
  signal blk00000001_sig000008ac : STD_LOGIC; 
  signal blk00000001_sig000008ab : STD_LOGIC; 
  signal blk00000001_sig000008aa : STD_LOGIC; 
  signal blk00000001_sig000008a9 : STD_LOGIC; 
  signal blk00000001_sig000008a8 : STD_LOGIC; 
  signal blk00000001_sig000008a7 : STD_LOGIC; 
  signal blk00000001_sig000008a6 : STD_LOGIC; 
  signal blk00000001_sig000008a5 : STD_LOGIC; 
  signal blk00000001_sig000008a4 : STD_LOGIC; 
  signal blk00000001_sig000008a3 : STD_LOGIC; 
  signal blk00000001_sig000008a2 : STD_LOGIC; 
  signal blk00000001_sig000008a1 : STD_LOGIC; 
  signal blk00000001_sig000008a0 : STD_LOGIC; 
  signal blk00000001_sig0000089f : STD_LOGIC; 
  signal blk00000001_sig0000089e : STD_LOGIC; 
  signal blk00000001_sig0000089d : STD_LOGIC; 
  signal blk00000001_sig0000089c : STD_LOGIC; 
  signal blk00000001_sig0000089b : STD_LOGIC; 
  signal blk00000001_sig0000089a : STD_LOGIC; 
  signal blk00000001_sig00000899 : STD_LOGIC; 
  signal blk00000001_sig00000898 : STD_LOGIC; 
  signal blk00000001_sig00000897 : STD_LOGIC; 
  signal blk00000001_sig00000896 : STD_LOGIC; 
  signal blk00000001_sig00000895 : STD_LOGIC; 
  signal blk00000001_sig00000894 : STD_LOGIC; 
  signal blk00000001_sig00000893 : STD_LOGIC; 
  signal blk00000001_sig00000892 : STD_LOGIC; 
  signal blk00000001_sig00000891 : STD_LOGIC; 
  signal blk00000001_sig00000890 : STD_LOGIC; 
  signal blk00000001_sig0000088f : STD_LOGIC; 
  signal blk00000001_sig0000088e : STD_LOGIC; 
  signal blk00000001_sig0000088d : STD_LOGIC; 
  signal blk00000001_sig0000088c : STD_LOGIC; 
  signal blk00000001_sig0000088b : STD_LOGIC; 
  signal blk00000001_sig0000088a : STD_LOGIC; 
  signal blk00000001_sig00000889 : STD_LOGIC; 
  signal blk00000001_sig00000888 : STD_LOGIC; 
  signal blk00000001_sig00000887 : STD_LOGIC; 
  signal blk00000001_sig00000886 : STD_LOGIC; 
  signal blk00000001_sig00000885 : STD_LOGIC; 
  signal blk00000001_sig00000884 : STD_LOGIC; 
  signal blk00000001_sig00000883 : STD_LOGIC; 
  signal blk00000001_sig00000882 : STD_LOGIC; 
  signal blk00000001_sig00000881 : STD_LOGIC; 
  signal blk00000001_sig00000880 : STD_LOGIC; 
  signal blk00000001_sig0000087f : STD_LOGIC; 
  signal blk00000001_sig0000087e : STD_LOGIC; 
  signal blk00000001_sig0000087d : STD_LOGIC; 
  signal blk00000001_sig0000087c : STD_LOGIC; 
  signal blk00000001_sig0000087b : STD_LOGIC; 
  signal blk00000001_sig0000087a : STD_LOGIC; 
  signal blk00000001_sig00000879 : STD_LOGIC; 
  signal blk00000001_sig00000878 : STD_LOGIC; 
  signal blk00000001_sig00000877 : STD_LOGIC; 
  signal blk00000001_sig00000876 : STD_LOGIC; 
  signal blk00000001_sig00000875 : STD_LOGIC; 
  signal blk00000001_sig00000874 : STD_LOGIC; 
  signal blk00000001_sig00000873 : STD_LOGIC; 
  signal blk00000001_sig00000872 : STD_LOGIC; 
  signal blk00000001_sig00000871 : STD_LOGIC; 
  signal blk00000001_sig00000870 : STD_LOGIC; 
  signal blk00000001_sig0000086f : STD_LOGIC; 
  signal blk00000001_sig0000086e : STD_LOGIC; 
  signal blk00000001_sig0000086d : STD_LOGIC; 
  signal blk00000001_sig0000086c : STD_LOGIC; 
  signal blk00000001_sig0000086b : STD_LOGIC; 
  signal blk00000001_sig0000086a : STD_LOGIC; 
  signal blk00000001_sig00000869 : STD_LOGIC; 
  signal blk00000001_sig00000868 : STD_LOGIC; 
  signal blk00000001_sig00000867 : STD_LOGIC; 
  signal blk00000001_sig00000866 : STD_LOGIC; 
  signal blk00000001_sig00000865 : STD_LOGIC; 
  signal blk00000001_sig00000864 : STD_LOGIC; 
  signal blk00000001_sig00000863 : STD_LOGIC; 
  signal blk00000001_sig00000862 : STD_LOGIC; 
  signal blk00000001_sig00000861 : STD_LOGIC; 
  signal blk00000001_sig00000860 : STD_LOGIC; 
  signal blk00000001_sig0000085f : STD_LOGIC; 
  signal blk00000001_sig0000085e : STD_LOGIC; 
  signal blk00000001_sig0000085d : STD_LOGIC; 
  signal blk00000001_sig0000085c : STD_LOGIC; 
  signal blk00000001_sig0000085b : STD_LOGIC; 
  signal blk00000001_sig0000085a : STD_LOGIC; 
  signal blk00000001_sig00000859 : STD_LOGIC; 
  signal blk00000001_sig00000858 : STD_LOGIC; 
  signal blk00000001_sig00000857 : STD_LOGIC; 
  signal blk00000001_sig00000856 : STD_LOGIC; 
  signal blk00000001_sig00000855 : STD_LOGIC; 
  signal blk00000001_sig00000854 : STD_LOGIC; 
  signal blk00000001_sig00000853 : STD_LOGIC; 
  signal blk00000001_sig00000852 : STD_LOGIC; 
  signal blk00000001_sig00000851 : STD_LOGIC; 
  signal blk00000001_sig00000850 : STD_LOGIC; 
  signal blk00000001_sig0000084f : STD_LOGIC; 
  signal blk00000001_sig0000084e : STD_LOGIC; 
  signal blk00000001_sig0000084d : STD_LOGIC; 
  signal blk00000001_sig0000084c : STD_LOGIC; 
  signal blk00000001_sig0000084b : STD_LOGIC; 
  signal blk00000001_sig0000084a : STD_LOGIC; 
  signal blk00000001_sig00000849 : STD_LOGIC; 
  signal blk00000001_sig00000848 : STD_LOGIC; 
  signal blk00000001_sig00000847 : STD_LOGIC; 
  signal blk00000001_sig00000846 : STD_LOGIC; 
  signal blk00000001_sig00000845 : STD_LOGIC; 
  signal blk00000001_sig00000844 : STD_LOGIC; 
  signal blk00000001_sig00000843 : STD_LOGIC; 
  signal blk00000001_sig00000842 : STD_LOGIC; 
  signal blk00000001_sig00000841 : STD_LOGIC; 
  signal blk00000001_sig00000840 : STD_LOGIC; 
  signal blk00000001_sig0000083f : STD_LOGIC; 
  signal blk00000001_sig0000083e : STD_LOGIC; 
  signal blk00000001_sig0000083d : STD_LOGIC; 
  signal blk00000001_sig0000083c : STD_LOGIC; 
  signal blk00000001_sig0000083b : STD_LOGIC; 
  signal blk00000001_sig0000083a : STD_LOGIC; 
  signal blk00000001_sig00000839 : STD_LOGIC; 
  signal blk00000001_sig00000838 : STD_LOGIC; 
  signal blk00000001_sig00000837 : STD_LOGIC; 
  signal blk00000001_sig00000836 : STD_LOGIC; 
  signal blk00000001_sig00000835 : STD_LOGIC; 
  signal blk00000001_sig00000834 : STD_LOGIC; 
  signal blk00000001_sig00000833 : STD_LOGIC; 
  signal blk00000001_sig00000832 : STD_LOGIC; 
  signal blk00000001_sig00000831 : STD_LOGIC; 
  signal blk00000001_sig00000830 : STD_LOGIC; 
  signal blk00000001_sig0000082f : STD_LOGIC; 
  signal blk00000001_sig0000082e : STD_LOGIC; 
  signal blk00000001_sig0000082d : STD_LOGIC; 
  signal blk00000001_sig0000082c : STD_LOGIC; 
  signal blk00000001_sig0000082b : STD_LOGIC; 
  signal blk00000001_sig0000082a : STD_LOGIC; 
  signal blk00000001_sig00000829 : STD_LOGIC; 
  signal blk00000001_sig00000828 : STD_LOGIC; 
  signal blk00000001_sig00000827 : STD_LOGIC; 
  signal blk00000001_sig00000826 : STD_LOGIC; 
  signal blk00000001_sig00000825 : STD_LOGIC; 
  signal blk00000001_sig00000824 : STD_LOGIC; 
  signal blk00000001_sig00000823 : STD_LOGIC; 
  signal blk00000001_sig00000822 : STD_LOGIC; 
  signal blk00000001_sig00000821 : STD_LOGIC; 
  signal blk00000001_sig00000820 : STD_LOGIC; 
  signal blk00000001_sig0000081f : STD_LOGIC; 
  signal blk00000001_sig0000081e : STD_LOGIC; 
  signal blk00000001_sig0000081d : STD_LOGIC; 
  signal blk00000001_sig0000081c : STD_LOGIC; 
  signal blk00000001_sig0000081b : STD_LOGIC; 
  signal blk00000001_sig0000081a : STD_LOGIC; 
  signal blk00000001_sig00000819 : STD_LOGIC; 
  signal blk00000001_sig00000818 : STD_LOGIC; 
  signal blk00000001_sig00000817 : STD_LOGIC; 
  signal blk00000001_sig00000816 : STD_LOGIC; 
  signal blk00000001_sig00000815 : STD_LOGIC; 
  signal blk00000001_sig00000814 : STD_LOGIC; 
  signal blk00000001_sig00000813 : STD_LOGIC; 
  signal blk00000001_sig00000812 : STD_LOGIC; 
  signal blk00000001_sig00000811 : STD_LOGIC; 
  signal blk00000001_sig00000810 : STD_LOGIC; 
  signal blk00000001_sig0000080f : STD_LOGIC; 
  signal blk00000001_sig0000080e : STD_LOGIC; 
  signal blk00000001_sig0000080d : STD_LOGIC; 
  signal blk00000001_sig0000080c : STD_LOGIC; 
  signal blk00000001_sig0000080b : STD_LOGIC; 
  signal blk00000001_sig0000080a : STD_LOGIC; 
  signal blk00000001_sig00000809 : STD_LOGIC; 
  signal blk00000001_sig00000808 : STD_LOGIC; 
  signal blk00000001_sig00000807 : STD_LOGIC; 
  signal blk00000001_sig00000806 : STD_LOGIC; 
  signal blk00000001_sig00000805 : STD_LOGIC; 
  signal blk00000001_sig00000804 : STD_LOGIC; 
  signal blk00000001_sig00000803 : STD_LOGIC; 
  signal blk00000001_sig00000802 : STD_LOGIC; 
  signal blk00000001_sig00000801 : STD_LOGIC; 
  signal blk00000001_sig00000800 : STD_LOGIC; 
  signal blk00000001_sig000007ff : STD_LOGIC; 
  signal blk00000001_sig000007fe : STD_LOGIC; 
  signal blk00000001_sig000007fd : STD_LOGIC; 
  signal blk00000001_sig000007fc : STD_LOGIC; 
  signal blk00000001_sig000007fb : STD_LOGIC; 
  signal blk00000001_sig000007fa : STD_LOGIC; 
  signal blk00000001_sig000007f9 : STD_LOGIC; 
  signal blk00000001_sig000007f8 : STD_LOGIC; 
  signal blk00000001_sig000007f7 : STD_LOGIC; 
  signal blk00000001_sig000007f6 : STD_LOGIC; 
  signal blk00000001_sig000007f5 : STD_LOGIC; 
  signal blk00000001_sig000007f4 : STD_LOGIC; 
  signal blk00000001_sig000007f3 : STD_LOGIC; 
  signal blk00000001_sig000007f2 : STD_LOGIC; 
  signal blk00000001_sig000007f1 : STD_LOGIC; 
  signal blk00000001_sig000007f0 : STD_LOGIC; 
  signal blk00000001_sig000007ef : STD_LOGIC; 
  signal blk00000001_sig000007ee : STD_LOGIC; 
  signal blk00000001_sig000007ed : STD_LOGIC; 
  signal blk00000001_sig000007ec : STD_LOGIC; 
  signal blk00000001_sig000007eb : STD_LOGIC; 
  signal blk00000001_sig000007ea : STD_LOGIC; 
  signal blk00000001_sig000007e9 : STD_LOGIC; 
  signal blk00000001_sig000007e8 : STD_LOGIC; 
  signal blk00000001_sig000007e7 : STD_LOGIC; 
  signal blk00000001_sig000007e6 : STD_LOGIC; 
  signal blk00000001_sig000007e5 : STD_LOGIC; 
  signal blk00000001_sig000007e4 : STD_LOGIC; 
  signal blk00000001_sig000007e3 : STD_LOGIC; 
  signal blk00000001_sig000007e2 : STD_LOGIC; 
  signal blk00000001_sig000007e1 : STD_LOGIC; 
  signal blk00000001_sig000007e0 : STD_LOGIC; 
  signal blk00000001_sig000007df : STD_LOGIC; 
  signal blk00000001_sig000007de : STD_LOGIC; 
  signal blk00000001_sig000007dd : STD_LOGIC; 
  signal blk00000001_sig000007dc : STD_LOGIC; 
  signal blk00000001_sig000007db : STD_LOGIC; 
  signal blk00000001_sig000007da : STD_LOGIC; 
  signal blk00000001_sig000007d9 : STD_LOGIC; 
  signal blk00000001_sig000007d8 : STD_LOGIC; 
  signal blk00000001_sig000007d7 : STD_LOGIC; 
  signal blk00000001_sig000007d6 : STD_LOGIC; 
  signal blk00000001_sig000007d5 : STD_LOGIC; 
  signal blk00000001_sig000007d4 : STD_LOGIC; 
  signal blk00000001_sig000007d3 : STD_LOGIC; 
  signal blk00000001_sig000007d2 : STD_LOGIC; 
  signal blk00000001_sig000007d1 : STD_LOGIC; 
  signal blk00000001_sig000007d0 : STD_LOGIC; 
  signal blk00000001_sig000007cf : STD_LOGIC; 
  signal blk00000001_sig000007ce : STD_LOGIC; 
  signal blk00000001_sig000007cd : STD_LOGIC; 
  signal blk00000001_sig000007cc : STD_LOGIC; 
  signal blk00000001_sig000007cb : STD_LOGIC; 
  signal blk00000001_sig000007ca : STD_LOGIC; 
  signal blk00000001_sig000007c9 : STD_LOGIC; 
  signal blk00000001_sig000007c8 : STD_LOGIC; 
  signal blk00000001_sig000007c7 : STD_LOGIC; 
  signal blk00000001_sig000007c6 : STD_LOGIC; 
  signal blk00000001_sig000007c5 : STD_LOGIC; 
  signal blk00000001_sig000007c4 : STD_LOGIC; 
  signal blk00000001_sig000007c3 : STD_LOGIC; 
  signal blk00000001_sig000007c2 : STD_LOGIC; 
  signal blk00000001_sig000007c1 : STD_LOGIC; 
  signal blk00000001_sig000007c0 : STD_LOGIC; 
  signal blk00000001_sig000007bf : STD_LOGIC; 
  signal blk00000001_sig000007be : STD_LOGIC; 
  signal blk00000001_sig000007bd : STD_LOGIC; 
  signal blk00000001_sig000007bc : STD_LOGIC; 
  signal blk00000001_sig000007bb : STD_LOGIC; 
  signal blk00000001_sig000007ba : STD_LOGIC; 
  signal blk00000001_sig000007b9 : STD_LOGIC; 
  signal blk00000001_sig000007b8 : STD_LOGIC; 
  signal blk00000001_sig000007b7 : STD_LOGIC; 
  signal blk00000001_sig000007b6 : STD_LOGIC; 
  signal blk00000001_sig000007b5 : STD_LOGIC; 
  signal blk00000001_sig000007b4 : STD_LOGIC; 
  signal blk00000001_sig000007b3 : STD_LOGIC; 
  signal blk00000001_sig000007b2 : STD_LOGIC; 
  signal blk00000001_sig000007b1 : STD_LOGIC; 
  signal blk00000001_sig000007b0 : STD_LOGIC; 
  signal blk00000001_sig000007af : STD_LOGIC; 
  signal blk00000001_sig000007ae : STD_LOGIC; 
  signal blk00000001_sig000007ad : STD_LOGIC; 
  signal blk00000001_sig000007ac : STD_LOGIC; 
  signal blk00000001_sig000007ab : STD_LOGIC; 
  signal blk00000001_sig000007aa : STD_LOGIC; 
  signal blk00000001_sig000007a9 : STD_LOGIC; 
  signal blk00000001_sig000007a8 : STD_LOGIC; 
  signal blk00000001_sig000007a7 : STD_LOGIC; 
  signal blk00000001_sig000007a6 : STD_LOGIC; 
  signal blk00000001_sig000007a5 : STD_LOGIC; 
  signal blk00000001_sig000007a4 : STD_LOGIC; 
  signal blk00000001_sig000007a3 : STD_LOGIC; 
  signal blk00000001_sig000007a2 : STD_LOGIC; 
  signal blk00000001_sig000007a1 : STD_LOGIC; 
  signal blk00000001_sig000007a0 : STD_LOGIC; 
  signal blk00000001_sig0000079f : STD_LOGIC; 
  signal blk00000001_sig0000079e : STD_LOGIC; 
  signal blk00000001_sig0000079d : STD_LOGIC; 
  signal blk00000001_sig0000079c : STD_LOGIC; 
  signal blk00000001_sig0000079b : STD_LOGIC; 
  signal blk00000001_sig0000079a : STD_LOGIC; 
  signal blk00000001_sig00000799 : STD_LOGIC; 
  signal blk00000001_sig00000798 : STD_LOGIC; 
  signal blk00000001_sig00000797 : STD_LOGIC; 
  signal blk00000001_sig00000796 : STD_LOGIC; 
  signal blk00000001_sig00000795 : STD_LOGIC; 
  signal blk00000001_sig00000794 : STD_LOGIC; 
  signal blk00000001_sig00000793 : STD_LOGIC; 
  signal blk00000001_sig00000792 : STD_LOGIC; 
  signal blk00000001_sig00000791 : STD_LOGIC; 
  signal blk00000001_sig00000790 : STD_LOGIC; 
  signal blk00000001_sig0000078f : STD_LOGIC; 
  signal blk00000001_sig0000078e : STD_LOGIC; 
  signal blk00000001_sig0000078d : STD_LOGIC; 
  signal blk00000001_sig0000078c : STD_LOGIC; 
  signal blk00000001_sig0000078b : STD_LOGIC; 
  signal blk00000001_sig0000078a : STD_LOGIC; 
  signal blk00000001_sig00000789 : STD_LOGIC; 
  signal blk00000001_sig00000788 : STD_LOGIC; 
  signal blk00000001_sig00000787 : STD_LOGIC; 
  signal blk00000001_sig00000786 : STD_LOGIC; 
  signal blk00000001_sig00000785 : STD_LOGIC; 
  signal blk00000001_sig00000784 : STD_LOGIC; 
  signal blk00000001_sig00000783 : STD_LOGIC; 
  signal blk00000001_sig00000782 : STD_LOGIC; 
  signal blk00000001_sig00000781 : STD_LOGIC; 
  signal blk00000001_sig00000780 : STD_LOGIC; 
  signal blk00000001_sig0000077f : STD_LOGIC; 
  signal blk00000001_sig0000077e : STD_LOGIC; 
  signal blk00000001_sig0000077d : STD_LOGIC; 
  signal blk00000001_sig0000077c : STD_LOGIC; 
  signal blk00000001_sig0000077b : STD_LOGIC; 
  signal blk00000001_sig0000077a : STD_LOGIC; 
  signal blk00000001_sig00000779 : STD_LOGIC; 
  signal blk00000001_sig00000778 : STD_LOGIC; 
  signal blk00000001_sig00000777 : STD_LOGIC; 
  signal blk00000001_sig00000776 : STD_LOGIC; 
  signal blk00000001_sig00000775 : STD_LOGIC; 
  signal blk00000001_sig00000774 : STD_LOGIC; 
  signal blk00000001_sig00000773 : STD_LOGIC; 
  signal blk00000001_sig00000772 : STD_LOGIC; 
  signal blk00000001_sig00000771 : STD_LOGIC; 
  signal blk00000001_sig00000770 : STD_LOGIC; 
  signal blk00000001_sig0000076f : STD_LOGIC; 
  signal blk00000001_sig0000076e : STD_LOGIC; 
  signal blk00000001_sig0000076d : STD_LOGIC; 
  signal blk00000001_sig0000076c : STD_LOGIC; 
  signal blk00000001_sig0000076b : STD_LOGIC; 
  signal blk00000001_sig0000076a : STD_LOGIC; 
  signal blk00000001_sig00000769 : STD_LOGIC; 
  signal blk00000001_sig00000768 : STD_LOGIC; 
  signal blk00000001_sig00000767 : STD_LOGIC; 
  signal blk00000001_sig00000766 : STD_LOGIC; 
  signal blk00000001_sig00000765 : STD_LOGIC; 
  signal blk00000001_sig00000764 : STD_LOGIC; 
  signal blk00000001_sig00000763 : STD_LOGIC; 
  signal blk00000001_sig00000762 : STD_LOGIC; 
  signal blk00000001_sig00000761 : STD_LOGIC; 
  signal blk00000001_sig00000760 : STD_LOGIC; 
  signal blk00000001_sig0000075f : STD_LOGIC; 
  signal blk00000001_sig0000075e : STD_LOGIC; 
  signal blk00000001_sig0000075d : STD_LOGIC; 
  signal blk00000001_sig0000075c : STD_LOGIC; 
  signal blk00000001_sig0000075b : STD_LOGIC; 
  signal blk00000001_sig0000075a : STD_LOGIC; 
  signal blk00000001_sig00000759 : STD_LOGIC; 
  signal blk00000001_sig00000758 : STD_LOGIC; 
  signal blk00000001_sig00000757 : STD_LOGIC; 
  signal blk00000001_sig00000756 : STD_LOGIC; 
  signal blk00000001_sig00000755 : STD_LOGIC; 
  signal blk00000001_sig00000754 : STD_LOGIC; 
  signal blk00000001_sig00000753 : STD_LOGIC; 
  signal blk00000001_sig00000752 : STD_LOGIC; 
  signal blk00000001_sig00000751 : STD_LOGIC; 
  signal blk00000001_sig00000750 : STD_LOGIC; 
  signal blk00000001_sig0000074f : STD_LOGIC; 
  signal blk00000001_sig0000074e : STD_LOGIC; 
  signal blk00000001_sig0000074d : STD_LOGIC; 
  signal blk00000001_sig0000074c : STD_LOGIC; 
  signal blk00000001_sig0000074b : STD_LOGIC; 
  signal blk00000001_sig0000074a : STD_LOGIC; 
  signal blk00000001_sig00000749 : STD_LOGIC; 
  signal blk00000001_sig00000748 : STD_LOGIC; 
  signal blk00000001_sig00000747 : STD_LOGIC; 
  signal blk00000001_sig00000746 : STD_LOGIC; 
  signal blk00000001_sig00000745 : STD_LOGIC; 
  signal blk00000001_sig00000744 : STD_LOGIC; 
  signal blk00000001_sig00000743 : STD_LOGIC; 
  signal blk00000001_sig00000742 : STD_LOGIC; 
  signal blk00000001_sig00000741 : STD_LOGIC; 
  signal blk00000001_sig00000740 : STD_LOGIC; 
  signal blk00000001_sig0000073f : STD_LOGIC; 
  signal blk00000001_sig0000073e : STD_LOGIC; 
  signal blk00000001_sig0000073d : STD_LOGIC; 
  signal blk00000001_sig0000073c : STD_LOGIC; 
  signal blk00000001_sig0000073b : STD_LOGIC; 
  signal blk00000001_sig0000073a : STD_LOGIC; 
  signal blk00000001_sig00000739 : STD_LOGIC; 
  signal blk00000001_sig00000738 : STD_LOGIC; 
  signal blk00000001_sig00000737 : STD_LOGIC; 
  signal blk00000001_sig00000736 : STD_LOGIC; 
  signal blk00000001_sig00000735 : STD_LOGIC; 
  signal blk00000001_sig00000734 : STD_LOGIC; 
  signal blk00000001_sig00000733 : STD_LOGIC; 
  signal blk00000001_sig00000732 : STD_LOGIC; 
  signal blk00000001_sig00000731 : STD_LOGIC; 
  signal blk00000001_sig00000730 : STD_LOGIC; 
  signal blk00000001_sig0000072f : STD_LOGIC; 
  signal blk00000001_sig0000072e : STD_LOGIC; 
  signal blk00000001_sig0000072d : STD_LOGIC; 
  signal blk00000001_sig0000072c : STD_LOGIC; 
  signal blk00000001_sig0000072b : STD_LOGIC; 
  signal blk00000001_sig0000072a : STD_LOGIC; 
  signal blk00000001_sig00000729 : STD_LOGIC; 
  signal blk00000001_sig00000728 : STD_LOGIC; 
  signal blk00000001_sig00000727 : STD_LOGIC; 
  signal blk00000001_sig00000726 : STD_LOGIC; 
  signal blk00000001_sig00000725 : STD_LOGIC; 
  signal blk00000001_sig00000724 : STD_LOGIC; 
  signal blk00000001_sig00000723 : STD_LOGIC; 
  signal blk00000001_sig00000722 : STD_LOGIC; 
  signal blk00000001_sig00000721 : STD_LOGIC; 
  signal blk00000001_sig00000720 : STD_LOGIC; 
  signal blk00000001_sig0000071f : STD_LOGIC; 
  signal blk00000001_sig0000071e : STD_LOGIC; 
  signal blk00000001_sig0000071d : STD_LOGIC; 
  signal blk00000001_sig0000071c : STD_LOGIC; 
  signal blk00000001_sig0000071b : STD_LOGIC; 
  signal blk00000001_sig0000071a : STD_LOGIC; 
  signal blk00000001_sig00000719 : STD_LOGIC; 
  signal blk00000001_sig00000718 : STD_LOGIC; 
  signal blk00000001_sig00000717 : STD_LOGIC; 
  signal blk00000001_sig00000716 : STD_LOGIC; 
  signal blk00000001_sig00000715 : STD_LOGIC; 
  signal blk00000001_sig00000714 : STD_LOGIC; 
  signal blk00000001_sig00000713 : STD_LOGIC; 
  signal blk00000001_sig00000712 : STD_LOGIC; 
  signal blk00000001_sig00000711 : STD_LOGIC; 
  signal blk00000001_sig00000710 : STD_LOGIC; 
  signal blk00000001_sig0000070f : STD_LOGIC; 
  signal blk00000001_sig0000070e : STD_LOGIC; 
  signal blk00000001_sig0000070d : STD_LOGIC; 
  signal blk00000001_sig0000070c : STD_LOGIC; 
  signal blk00000001_sig0000070b : STD_LOGIC; 
  signal blk00000001_sig0000070a : STD_LOGIC; 
  signal blk00000001_sig00000709 : STD_LOGIC; 
  signal blk00000001_sig00000708 : STD_LOGIC; 
  signal blk00000001_sig00000707 : STD_LOGIC; 
  signal blk00000001_sig00000706 : STD_LOGIC; 
  signal blk00000001_sig00000705 : STD_LOGIC; 
  signal blk00000001_sig00000704 : STD_LOGIC; 
  signal blk00000001_sig00000703 : STD_LOGIC; 
  signal blk00000001_sig00000702 : STD_LOGIC; 
  signal blk00000001_sig00000701 : STD_LOGIC; 
  signal blk00000001_sig00000700 : STD_LOGIC; 
  signal blk00000001_sig000006ff : STD_LOGIC; 
  signal blk00000001_sig000006fe : STD_LOGIC; 
  signal blk00000001_sig000006fd : STD_LOGIC; 
  signal blk00000001_sig000006fc : STD_LOGIC; 
  signal blk00000001_sig000006fb : STD_LOGIC; 
  signal blk00000001_sig000006fa : STD_LOGIC; 
  signal blk00000001_sig000006f9 : STD_LOGIC; 
  signal blk00000001_sig000006f8 : STD_LOGIC; 
  signal blk00000001_sig000006f7 : STD_LOGIC; 
  signal blk00000001_sig000006f6 : STD_LOGIC; 
  signal blk00000001_sig000006f5 : STD_LOGIC; 
  signal blk00000001_sig000006f4 : STD_LOGIC; 
  signal blk00000001_sig000006f3 : STD_LOGIC; 
  signal blk00000001_sig000006f2 : STD_LOGIC; 
  signal blk00000001_sig000006f1 : STD_LOGIC; 
  signal blk00000001_sig000006f0 : STD_LOGIC; 
  signal blk00000001_sig000006ef : STD_LOGIC; 
  signal blk00000001_sig000006ee : STD_LOGIC; 
  signal blk00000001_sig000006ed : STD_LOGIC; 
  signal blk00000001_sig000006ec : STD_LOGIC; 
  signal blk00000001_sig000006eb : STD_LOGIC; 
  signal blk00000001_sig000006ea : STD_LOGIC; 
  signal blk00000001_sig000006e9 : STD_LOGIC; 
  signal blk00000001_sig000006e8 : STD_LOGIC; 
  signal blk00000001_sig000006e7 : STD_LOGIC; 
  signal blk00000001_sig000006e6 : STD_LOGIC; 
  signal blk00000001_sig000006e5 : STD_LOGIC; 
  signal blk00000001_sig000006e4 : STD_LOGIC; 
  signal blk00000001_sig000006e3 : STD_LOGIC; 
  signal blk00000001_sig000006e2 : STD_LOGIC; 
  signal blk00000001_sig000006e1 : STD_LOGIC; 
  signal blk00000001_sig000006e0 : STD_LOGIC; 
  signal blk00000001_sig000006df : STD_LOGIC; 
  signal blk00000001_sig000006de : STD_LOGIC; 
  signal blk00000001_sig000006dd : STD_LOGIC; 
  signal blk00000001_sig000006dc : STD_LOGIC; 
  signal blk00000001_sig000006db : STD_LOGIC; 
  signal blk00000001_sig000006da : STD_LOGIC; 
  signal blk00000001_sig000006d9 : STD_LOGIC; 
  signal blk00000001_sig000006d8 : STD_LOGIC; 
  signal blk00000001_sig000006d7 : STD_LOGIC; 
  signal blk00000001_sig000006d6 : STD_LOGIC; 
  signal blk00000001_sig000006d5 : STD_LOGIC; 
  signal blk00000001_sig000006d4 : STD_LOGIC; 
  signal blk00000001_sig000006d3 : STD_LOGIC; 
  signal blk00000001_sig000006d2 : STD_LOGIC; 
  signal blk00000001_sig000006d1 : STD_LOGIC; 
  signal blk00000001_sig000006d0 : STD_LOGIC; 
  signal blk00000001_sig000006cf : STD_LOGIC; 
  signal blk00000001_sig000006ce : STD_LOGIC; 
  signal blk00000001_sig000006cd : STD_LOGIC; 
  signal blk00000001_sig000006cc : STD_LOGIC; 
  signal blk00000001_sig000006cb : STD_LOGIC; 
  signal blk00000001_sig000006ca : STD_LOGIC; 
  signal blk00000001_sig000006c9 : STD_LOGIC; 
  signal blk00000001_sig000006c8 : STD_LOGIC; 
  signal blk00000001_sig000006c7 : STD_LOGIC; 
  signal blk00000001_sig000006c6 : STD_LOGIC; 
  signal blk00000001_sig000006c5 : STD_LOGIC; 
  signal blk00000001_sig000006c4 : STD_LOGIC; 
  signal blk00000001_sig000006c3 : STD_LOGIC; 
  signal blk00000001_sig000006c2 : STD_LOGIC; 
  signal blk00000001_sig000006c1 : STD_LOGIC; 
  signal blk00000001_sig000006c0 : STD_LOGIC; 
  signal blk00000001_sig000006bf : STD_LOGIC; 
  signal blk00000001_sig000006be : STD_LOGIC; 
  signal blk00000001_sig000006bd : STD_LOGIC; 
  signal blk00000001_sig000006bc : STD_LOGIC; 
  signal blk00000001_sig000006bb : STD_LOGIC; 
  signal blk00000001_sig000006ba : STD_LOGIC; 
  signal blk00000001_sig000006b9 : STD_LOGIC; 
  signal blk00000001_sig000006b8 : STD_LOGIC; 
  signal blk00000001_sig000006b7 : STD_LOGIC; 
  signal blk00000001_sig000006b6 : STD_LOGIC; 
  signal blk00000001_sig000006b5 : STD_LOGIC; 
  signal blk00000001_sig000006b4 : STD_LOGIC; 
  signal blk00000001_sig000006b3 : STD_LOGIC; 
  signal blk00000001_sig000006b2 : STD_LOGIC; 
  signal blk00000001_sig000006b1 : STD_LOGIC; 
  signal blk00000001_sig000006b0 : STD_LOGIC; 
  signal blk00000001_sig000006af : STD_LOGIC; 
  signal blk00000001_sig000006ae : STD_LOGIC; 
  signal blk00000001_sig000006ad : STD_LOGIC; 
  signal blk00000001_sig000006ac : STD_LOGIC; 
  signal blk00000001_sig000006ab : STD_LOGIC; 
  signal blk00000001_sig000006aa : STD_LOGIC; 
  signal blk00000001_sig000006a9 : STD_LOGIC; 
  signal blk00000001_sig000006a8 : STD_LOGIC; 
  signal blk00000001_sig000006a7 : STD_LOGIC; 
  signal blk00000001_sig000006a6 : STD_LOGIC; 
  signal blk00000001_sig000006a5 : STD_LOGIC; 
  signal blk00000001_sig000006a4 : STD_LOGIC; 
  signal blk00000001_sig000006a3 : STD_LOGIC; 
  signal blk00000001_sig000006a2 : STD_LOGIC; 
  signal blk00000001_sig000006a1 : STD_LOGIC; 
  signal blk00000001_sig000006a0 : STD_LOGIC; 
  signal blk00000001_sig0000069f : STD_LOGIC; 
  signal blk00000001_sig0000069e : STD_LOGIC; 
  signal blk00000001_sig0000069d : STD_LOGIC; 
  signal blk00000001_sig0000069c : STD_LOGIC; 
  signal blk00000001_sig0000069b : STD_LOGIC; 
  signal blk00000001_sig0000069a : STD_LOGIC; 
  signal blk00000001_sig00000699 : STD_LOGIC; 
  signal blk00000001_sig00000698 : STD_LOGIC; 
  signal blk00000001_sig00000697 : STD_LOGIC; 
  signal blk00000001_sig00000696 : STD_LOGIC; 
  signal blk00000001_sig00000695 : STD_LOGIC; 
  signal blk00000001_sig00000694 : STD_LOGIC; 
  signal blk00000001_sig00000693 : STD_LOGIC; 
  signal blk00000001_sig00000692 : STD_LOGIC; 
  signal blk00000001_sig00000691 : STD_LOGIC; 
  signal blk00000001_sig00000690 : STD_LOGIC; 
  signal blk00000001_sig0000068f : STD_LOGIC; 
  signal blk00000001_sig0000068e : STD_LOGIC; 
  signal blk00000001_sig0000068d : STD_LOGIC; 
  signal blk00000001_sig0000068c : STD_LOGIC; 
  signal blk00000001_sig0000068b : STD_LOGIC; 
  signal blk00000001_sig0000068a : STD_LOGIC; 
  signal blk00000001_sig00000689 : STD_LOGIC; 
  signal blk00000001_sig00000688 : STD_LOGIC; 
  signal blk00000001_sig00000687 : STD_LOGIC; 
  signal blk00000001_sig00000686 : STD_LOGIC; 
  signal blk00000001_sig00000685 : STD_LOGIC; 
  signal blk00000001_sig00000684 : STD_LOGIC; 
  signal blk00000001_sig00000683 : STD_LOGIC; 
  signal blk00000001_sig00000682 : STD_LOGIC; 
  signal blk00000001_sig00000681 : STD_LOGIC; 
  signal blk00000001_sig00000680 : STD_LOGIC; 
  signal blk00000001_sig0000067f : STD_LOGIC; 
  signal blk00000001_sig0000067e : STD_LOGIC; 
  signal blk00000001_sig0000067d : STD_LOGIC; 
  signal blk00000001_sig0000067c : STD_LOGIC; 
  signal blk00000001_sig0000067b : STD_LOGIC; 
  signal blk00000001_sig0000067a : STD_LOGIC; 
  signal blk00000001_sig00000679 : STD_LOGIC; 
  signal blk00000001_sig00000678 : STD_LOGIC; 
  signal blk00000001_sig00000677 : STD_LOGIC; 
  signal blk00000001_sig00000676 : STD_LOGIC; 
  signal blk00000001_sig00000675 : STD_LOGIC; 
  signal blk00000001_sig00000674 : STD_LOGIC; 
  signal blk00000001_sig00000673 : STD_LOGIC; 
  signal blk00000001_sig00000672 : STD_LOGIC; 
  signal blk00000001_sig00000671 : STD_LOGIC; 
  signal blk00000001_sig00000670 : STD_LOGIC; 
  signal blk00000001_sig0000066f : STD_LOGIC; 
  signal blk00000001_sig0000066e : STD_LOGIC; 
  signal blk00000001_sig0000066d : STD_LOGIC; 
  signal blk00000001_sig0000066c : STD_LOGIC; 
  signal blk00000001_sig0000066b : STD_LOGIC; 
  signal blk00000001_sig0000066a : STD_LOGIC; 
  signal blk00000001_sig00000669 : STD_LOGIC; 
  signal blk00000001_sig00000668 : STD_LOGIC; 
  signal blk00000001_sig00000667 : STD_LOGIC; 
  signal blk00000001_sig00000666 : STD_LOGIC; 
  signal blk00000001_sig00000665 : STD_LOGIC; 
  signal blk00000001_sig00000664 : STD_LOGIC; 
  signal blk00000001_sig00000663 : STD_LOGIC; 
  signal blk00000001_sig00000662 : STD_LOGIC; 
  signal blk00000001_sig00000661 : STD_LOGIC; 
  signal blk00000001_sig00000660 : STD_LOGIC; 
  signal blk00000001_sig0000065f : STD_LOGIC; 
  signal blk00000001_sig0000065e : STD_LOGIC; 
  signal blk00000001_sig0000065d : STD_LOGIC; 
  signal blk00000001_sig0000065c : STD_LOGIC; 
  signal blk00000001_sig0000065b : STD_LOGIC; 
  signal blk00000001_sig0000065a : STD_LOGIC; 
  signal blk00000001_sig00000659 : STD_LOGIC; 
  signal blk00000001_sig00000658 : STD_LOGIC; 
  signal blk00000001_sig00000657 : STD_LOGIC; 
  signal blk00000001_sig00000656 : STD_LOGIC; 
  signal blk00000001_sig00000655 : STD_LOGIC; 
  signal blk00000001_sig00000654 : STD_LOGIC; 
  signal blk00000001_sig00000653 : STD_LOGIC; 
  signal blk00000001_sig00000652 : STD_LOGIC; 
  signal blk00000001_sig00000651 : STD_LOGIC; 
  signal blk00000001_sig00000650 : STD_LOGIC; 
  signal blk00000001_sig0000064f : STD_LOGIC; 
  signal blk00000001_sig0000064e : STD_LOGIC; 
  signal blk00000001_sig0000064d : STD_LOGIC; 
  signal blk00000001_sig0000064c : STD_LOGIC; 
  signal blk00000001_sig0000064b : STD_LOGIC; 
  signal blk00000001_sig0000064a : STD_LOGIC; 
  signal blk00000001_sig00000649 : STD_LOGIC; 
  signal blk00000001_sig00000648 : STD_LOGIC; 
  signal blk00000001_sig00000647 : STD_LOGIC; 
  signal blk00000001_sig00000646 : STD_LOGIC; 
  signal blk00000001_sig00000645 : STD_LOGIC; 
  signal blk00000001_sig00000644 : STD_LOGIC; 
  signal blk00000001_sig00000643 : STD_LOGIC; 
  signal blk00000001_sig00000642 : STD_LOGIC; 
  signal blk00000001_sig00000641 : STD_LOGIC; 
  signal blk00000001_sig00000640 : STD_LOGIC; 
  signal blk00000001_sig0000063f : STD_LOGIC; 
  signal blk00000001_sig0000063e : STD_LOGIC; 
  signal blk00000001_sig0000063d : STD_LOGIC; 
  signal blk00000001_sig0000063c : STD_LOGIC; 
  signal blk00000001_sig0000063b : STD_LOGIC; 
  signal blk00000001_sig0000063a : STD_LOGIC; 
  signal blk00000001_sig00000639 : STD_LOGIC; 
  signal blk00000001_sig00000638 : STD_LOGIC; 
  signal blk00000001_sig00000637 : STD_LOGIC; 
  signal blk00000001_sig00000636 : STD_LOGIC; 
  signal blk00000001_sig00000635 : STD_LOGIC; 
  signal blk00000001_sig00000634 : STD_LOGIC; 
  signal blk00000001_sig00000633 : STD_LOGIC; 
  signal blk00000001_sig00000632 : STD_LOGIC; 
  signal blk00000001_sig00000631 : STD_LOGIC; 
  signal blk00000001_sig00000630 : STD_LOGIC; 
  signal blk00000001_sig0000062f : STD_LOGIC; 
  signal blk00000001_sig0000062e : STD_LOGIC; 
  signal blk00000001_sig0000062d : STD_LOGIC; 
  signal blk00000001_sig0000062c : STD_LOGIC; 
  signal blk00000001_sig0000062b : STD_LOGIC; 
  signal blk00000001_sig0000062a : STD_LOGIC; 
  signal blk00000001_sig00000629 : STD_LOGIC; 
  signal blk00000001_sig00000628 : STD_LOGIC; 
  signal blk00000001_sig00000627 : STD_LOGIC; 
  signal blk00000001_sig00000626 : STD_LOGIC; 
  signal blk00000001_sig00000625 : STD_LOGIC; 
  signal blk00000001_sig00000624 : STD_LOGIC; 
  signal blk00000001_sig00000623 : STD_LOGIC; 
  signal blk00000001_sig00000622 : STD_LOGIC; 
  signal blk00000001_sig00000621 : STD_LOGIC; 
  signal blk00000001_sig00000620 : STD_LOGIC; 
  signal blk00000001_sig0000061f : STD_LOGIC; 
  signal blk00000001_sig0000061e : STD_LOGIC; 
  signal blk00000001_sig0000061d : STD_LOGIC; 
  signal blk00000001_sig0000061c : STD_LOGIC; 
  signal blk00000001_sig0000061b : STD_LOGIC; 
  signal blk00000001_sig0000061a : STD_LOGIC; 
  signal blk00000001_sig00000619 : STD_LOGIC; 
  signal blk00000001_sig00000618 : STD_LOGIC; 
  signal blk00000001_sig00000617 : STD_LOGIC; 
  signal blk00000001_sig00000616 : STD_LOGIC; 
  signal blk00000001_sig00000615 : STD_LOGIC; 
  signal blk00000001_sig00000614 : STD_LOGIC; 
  signal blk00000001_sig00000613 : STD_LOGIC; 
  signal blk00000001_sig00000612 : STD_LOGIC; 
  signal blk00000001_sig00000611 : STD_LOGIC; 
  signal blk00000001_sig00000610 : STD_LOGIC; 
  signal blk00000001_sig0000060f : STD_LOGIC; 
  signal blk00000001_sig0000060e : STD_LOGIC; 
  signal blk00000001_sig0000060d : STD_LOGIC; 
  signal blk00000001_sig0000060c : STD_LOGIC; 
  signal blk00000001_sig0000060b : STD_LOGIC; 
  signal blk00000001_sig0000060a : STD_LOGIC; 
  signal blk00000001_sig00000609 : STD_LOGIC; 
  signal blk00000001_sig00000608 : STD_LOGIC; 
  signal blk00000001_sig00000607 : STD_LOGIC; 
  signal blk00000001_sig00000606 : STD_LOGIC; 
  signal blk00000001_sig00000605 : STD_LOGIC; 
  signal blk00000001_sig00000604 : STD_LOGIC; 
  signal blk00000001_sig00000603 : STD_LOGIC; 
  signal blk00000001_sig00000602 : STD_LOGIC; 
  signal blk00000001_sig00000601 : STD_LOGIC; 
  signal blk00000001_sig00000600 : STD_LOGIC; 
  signal blk00000001_sig000005ff : STD_LOGIC; 
  signal blk00000001_sig000005fe : STD_LOGIC; 
  signal blk00000001_sig000005fd : STD_LOGIC; 
  signal blk00000001_sig000005fc : STD_LOGIC; 
  signal blk00000001_sig000005fb : STD_LOGIC; 
  signal blk00000001_sig000005fa : STD_LOGIC; 
  signal blk00000001_sig000005f9 : STD_LOGIC; 
  signal blk00000001_sig000005f8 : STD_LOGIC; 
  signal blk00000001_sig000005f7 : STD_LOGIC; 
  signal blk00000001_sig000005f6 : STD_LOGIC; 
  signal blk00000001_sig000005f5 : STD_LOGIC; 
  signal blk00000001_sig000005f4 : STD_LOGIC; 
  signal blk00000001_sig000005f3 : STD_LOGIC; 
  signal blk00000001_sig000005f2 : STD_LOGIC; 
  signal blk00000001_sig000005f1 : STD_LOGIC; 
  signal blk00000001_sig000005f0 : STD_LOGIC; 
  signal blk00000001_sig000005ef : STD_LOGIC; 
  signal blk00000001_sig000005ee : STD_LOGIC; 
  signal blk00000001_sig000005ed : STD_LOGIC; 
  signal blk00000001_sig000005ec : STD_LOGIC; 
  signal blk00000001_sig000005eb : STD_LOGIC; 
  signal blk00000001_sig000005ea : STD_LOGIC; 
  signal blk00000001_sig000005e9 : STD_LOGIC; 
  signal blk00000001_sig000005e8 : STD_LOGIC; 
  signal blk00000001_sig000005e7 : STD_LOGIC; 
  signal blk00000001_sig000005e6 : STD_LOGIC; 
  signal blk00000001_sig000005e5 : STD_LOGIC; 
  signal blk00000001_sig000005e4 : STD_LOGIC; 
  signal blk00000001_sig000005e3 : STD_LOGIC; 
  signal blk00000001_sig000005e2 : STD_LOGIC; 
  signal blk00000001_sig000005e1 : STD_LOGIC; 
  signal blk00000001_sig000005e0 : STD_LOGIC; 
  signal blk00000001_sig000005df : STD_LOGIC; 
  signal blk00000001_sig000005de : STD_LOGIC; 
  signal blk00000001_sig000005dd : STD_LOGIC; 
  signal blk00000001_sig000005dc : STD_LOGIC; 
  signal blk00000001_sig000005db : STD_LOGIC; 
  signal blk00000001_sig000005da : STD_LOGIC; 
  signal blk00000001_sig000005d9 : STD_LOGIC; 
  signal blk00000001_sig000005d8 : STD_LOGIC; 
  signal blk00000001_sig000005d7 : STD_LOGIC; 
  signal blk00000001_sig000005d6 : STD_LOGIC; 
  signal blk00000001_sig000005d5 : STD_LOGIC; 
  signal blk00000001_sig000005d4 : STD_LOGIC; 
  signal blk00000001_sig000005d3 : STD_LOGIC; 
  signal blk00000001_sig000005d2 : STD_LOGIC; 
  signal blk00000001_sig000005d1 : STD_LOGIC; 
  signal blk00000001_sig000005d0 : STD_LOGIC; 
  signal blk00000001_sig000005cf : STD_LOGIC; 
  signal blk00000001_sig000005ce : STD_LOGIC; 
  signal blk00000001_sig000005cd : STD_LOGIC; 
  signal blk00000001_sig000005cc : STD_LOGIC; 
  signal blk00000001_sig000005cb : STD_LOGIC; 
  signal blk00000001_sig000005ca : STD_LOGIC; 
  signal blk00000001_sig000005c9 : STD_LOGIC; 
  signal blk00000001_sig000005c8 : STD_LOGIC; 
  signal blk00000001_sig000005c7 : STD_LOGIC; 
  signal blk00000001_sig000005c6 : STD_LOGIC; 
  signal blk00000001_sig000005c5 : STD_LOGIC; 
  signal blk00000001_sig000005c4 : STD_LOGIC; 
  signal blk00000001_sig000005c3 : STD_LOGIC; 
  signal blk00000001_sig000005c2 : STD_LOGIC; 
  signal blk00000001_sig000005c1 : STD_LOGIC; 
  signal blk00000001_sig000005c0 : STD_LOGIC; 
  signal blk00000001_sig000005bf : STD_LOGIC; 
  signal blk00000001_sig000005be : STD_LOGIC; 
  signal blk00000001_sig000005bd : STD_LOGIC; 
  signal blk00000001_sig000005bc : STD_LOGIC; 
  signal blk00000001_sig000005bb : STD_LOGIC; 
  signal blk00000001_sig000005ba : STD_LOGIC; 
  signal blk00000001_sig000005b9 : STD_LOGIC; 
  signal blk00000001_sig000005b8 : STD_LOGIC; 
  signal blk00000001_sig000005b7 : STD_LOGIC; 
  signal blk00000001_sig000005b6 : STD_LOGIC; 
  signal blk00000001_sig000005b5 : STD_LOGIC; 
  signal blk00000001_sig000005b4 : STD_LOGIC; 
  signal blk00000001_sig000005b3 : STD_LOGIC; 
  signal blk00000001_sig000005b2 : STD_LOGIC; 
  signal blk00000001_sig000005b1 : STD_LOGIC; 
  signal blk00000001_sig000005b0 : STD_LOGIC; 
  signal blk00000001_sig000005af : STD_LOGIC; 
  signal blk00000001_sig000005ae : STD_LOGIC; 
  signal blk00000001_sig000005ad : STD_LOGIC; 
  signal blk00000001_sig000005ac : STD_LOGIC; 
  signal blk00000001_sig000005ab : STD_LOGIC; 
  signal blk00000001_sig000005aa : STD_LOGIC; 
  signal blk00000001_sig000005a9 : STD_LOGIC; 
  signal blk00000001_sig000005a8 : STD_LOGIC; 
  signal blk00000001_sig000005a7 : STD_LOGIC; 
  signal blk00000001_sig000005a6 : STD_LOGIC; 
  signal blk00000001_sig000005a5 : STD_LOGIC; 
  signal blk00000001_sig000005a4 : STD_LOGIC; 
  signal blk00000001_sig000005a3 : STD_LOGIC; 
  signal blk00000001_sig000005a2 : STD_LOGIC; 
  signal blk00000001_sig000005a1 : STD_LOGIC; 
  signal blk00000001_sig000005a0 : STD_LOGIC; 
  signal blk00000001_sig0000059f : STD_LOGIC; 
  signal blk00000001_sig0000059e : STD_LOGIC; 
  signal blk00000001_sig0000059d : STD_LOGIC; 
  signal blk00000001_sig0000059c : STD_LOGIC; 
  signal blk00000001_sig0000059b : STD_LOGIC; 
  signal blk00000001_sig0000059a : STD_LOGIC; 
  signal blk00000001_sig00000599 : STD_LOGIC; 
  signal blk00000001_sig00000598 : STD_LOGIC; 
  signal blk00000001_sig00000597 : STD_LOGIC; 
  signal blk00000001_sig00000596 : STD_LOGIC; 
  signal blk00000001_sig00000595 : STD_LOGIC; 
  signal blk00000001_sig00000594 : STD_LOGIC; 
  signal blk00000001_sig00000593 : STD_LOGIC; 
  signal blk00000001_sig00000592 : STD_LOGIC; 
  signal blk00000001_sig00000591 : STD_LOGIC; 
  signal blk00000001_sig00000590 : STD_LOGIC; 
  signal blk00000001_sig0000058f : STD_LOGIC; 
  signal blk00000001_sig0000058e : STD_LOGIC; 
  signal blk00000001_sig0000058d : STD_LOGIC; 
  signal blk00000001_sig0000058c : STD_LOGIC; 
  signal blk00000001_sig0000058b : STD_LOGIC; 
  signal blk00000001_sig0000058a : STD_LOGIC; 
  signal blk00000001_sig00000589 : STD_LOGIC; 
  signal blk00000001_sig00000588 : STD_LOGIC; 
  signal blk00000001_sig00000587 : STD_LOGIC; 
  signal blk00000001_sig00000586 : STD_LOGIC; 
  signal blk00000001_sig00000585 : STD_LOGIC; 
  signal blk00000001_sig00000584 : STD_LOGIC; 
  signal blk00000001_sig00000583 : STD_LOGIC; 
  signal blk00000001_sig00000582 : STD_LOGIC; 
  signal blk00000001_sig00000581 : STD_LOGIC; 
  signal blk00000001_sig00000580 : STD_LOGIC; 
  signal blk00000001_sig0000057f : STD_LOGIC; 
  signal blk00000001_sig0000057e : STD_LOGIC; 
  signal blk00000001_sig0000057d : STD_LOGIC; 
  signal blk00000001_sig0000057c : STD_LOGIC; 
  signal blk00000001_sig0000057b : STD_LOGIC; 
  signal blk00000001_sig0000057a : STD_LOGIC; 
  signal blk00000001_sig00000579 : STD_LOGIC; 
  signal blk00000001_sig00000578 : STD_LOGIC; 
  signal blk00000001_sig00000577 : STD_LOGIC; 
  signal blk00000001_sig00000576 : STD_LOGIC; 
  signal blk00000001_sig00000575 : STD_LOGIC; 
  signal blk00000001_sig00000574 : STD_LOGIC; 
  signal blk00000001_sig00000573 : STD_LOGIC; 
  signal blk00000001_sig00000572 : STD_LOGIC; 
  signal blk00000001_sig00000571 : STD_LOGIC; 
  signal blk00000001_sig00000570 : STD_LOGIC; 
  signal blk00000001_sig0000056f : STD_LOGIC; 
  signal blk00000001_sig0000056e : STD_LOGIC; 
  signal blk00000001_sig0000056d : STD_LOGIC; 
  signal blk00000001_sig0000056c : STD_LOGIC; 
  signal blk00000001_sig0000056b : STD_LOGIC; 
  signal blk00000001_sig0000056a : STD_LOGIC; 
  signal blk00000001_sig00000569 : STD_LOGIC; 
  signal blk00000001_sig00000568 : STD_LOGIC; 
  signal blk00000001_sig00000567 : STD_LOGIC; 
  signal blk00000001_sig00000566 : STD_LOGIC; 
  signal blk00000001_sig00000565 : STD_LOGIC; 
  signal blk00000001_sig00000564 : STD_LOGIC; 
  signal blk00000001_sig00000563 : STD_LOGIC; 
  signal blk00000001_sig00000562 : STD_LOGIC; 
  signal blk00000001_sig00000561 : STD_LOGIC; 
  signal blk00000001_sig00000560 : STD_LOGIC; 
  signal blk00000001_sig0000055f : STD_LOGIC; 
  signal blk00000001_sig0000055e : STD_LOGIC; 
  signal blk00000001_sig0000055d : STD_LOGIC; 
  signal blk00000001_sig0000055c : STD_LOGIC; 
  signal blk00000001_sig0000055b : STD_LOGIC; 
  signal blk00000001_sig0000055a : STD_LOGIC; 
  signal blk00000001_sig00000559 : STD_LOGIC; 
  signal blk00000001_sig00000558 : STD_LOGIC; 
  signal blk00000001_sig00000557 : STD_LOGIC; 
  signal blk00000001_sig00000556 : STD_LOGIC; 
  signal blk00000001_sig00000555 : STD_LOGIC; 
  signal blk00000001_sig00000554 : STD_LOGIC; 
  signal blk00000001_sig00000553 : STD_LOGIC; 
  signal blk00000001_sig00000552 : STD_LOGIC; 
  signal blk00000001_sig00000551 : STD_LOGIC; 
  signal blk00000001_sig00000550 : STD_LOGIC; 
  signal blk00000001_sig0000054f : STD_LOGIC; 
  signal blk00000001_sig0000054e : STD_LOGIC; 
  signal blk00000001_sig0000054d : STD_LOGIC; 
  signal blk00000001_sig0000054c : STD_LOGIC; 
  signal blk00000001_sig0000054b : STD_LOGIC; 
  signal blk00000001_sig0000054a : STD_LOGIC; 
  signal blk00000001_sig00000549 : STD_LOGIC; 
  signal blk00000001_sig00000548 : STD_LOGIC; 
  signal blk00000001_sig00000547 : STD_LOGIC; 
  signal blk00000001_sig00000546 : STD_LOGIC; 
  signal blk00000001_sig00000545 : STD_LOGIC; 
  signal blk00000001_sig00000544 : STD_LOGIC; 
  signal blk00000001_sig00000543 : STD_LOGIC; 
  signal blk00000001_sig00000542 : STD_LOGIC; 
  signal blk00000001_sig00000541 : STD_LOGIC; 
  signal blk00000001_sig00000540 : STD_LOGIC; 
  signal blk00000001_sig0000053f : STD_LOGIC; 
  signal blk00000001_sig0000053e : STD_LOGIC; 
  signal blk00000001_sig0000053d : STD_LOGIC; 
  signal blk00000001_sig0000053c : STD_LOGIC; 
  signal blk00000001_sig0000053b : STD_LOGIC; 
  signal blk00000001_sig0000053a : STD_LOGIC; 
  signal blk00000001_sig00000539 : STD_LOGIC; 
  signal blk00000001_sig00000538 : STD_LOGIC; 
  signal blk00000001_sig00000537 : STD_LOGIC; 
  signal blk00000001_sig00000536 : STD_LOGIC; 
  signal blk00000001_sig00000535 : STD_LOGIC; 
  signal blk00000001_sig00000534 : STD_LOGIC; 
  signal blk00000001_sig00000533 : STD_LOGIC; 
  signal blk00000001_sig00000532 : STD_LOGIC; 
  signal blk00000001_sig00000531 : STD_LOGIC; 
  signal blk00000001_sig00000530 : STD_LOGIC; 
  signal blk00000001_sig0000052f : STD_LOGIC; 
  signal blk00000001_sig0000052e : STD_LOGIC; 
  signal blk00000001_sig0000052d : STD_LOGIC; 
  signal blk00000001_sig0000052c : STD_LOGIC; 
  signal blk00000001_sig0000052b : STD_LOGIC; 
  signal blk00000001_sig0000052a : STD_LOGIC; 
  signal blk00000001_sig00000529 : STD_LOGIC; 
  signal blk00000001_sig00000528 : STD_LOGIC; 
  signal blk00000001_sig00000527 : STD_LOGIC; 
  signal blk00000001_sig00000526 : STD_LOGIC; 
  signal blk00000001_sig00000525 : STD_LOGIC; 
  signal blk00000001_sig00000524 : STD_LOGIC; 
  signal blk00000001_sig00000523 : STD_LOGIC; 
  signal blk00000001_sig00000522 : STD_LOGIC; 
  signal blk00000001_sig00000521 : STD_LOGIC; 
  signal blk00000001_sig00000520 : STD_LOGIC; 
  signal blk00000001_sig0000051f : STD_LOGIC; 
  signal blk00000001_sig0000051e : STD_LOGIC; 
  signal blk00000001_sig0000051d : STD_LOGIC; 
  signal blk00000001_sig0000051c : STD_LOGIC; 
  signal blk00000001_sig0000051b : STD_LOGIC; 
  signal blk00000001_sig0000051a : STD_LOGIC; 
  signal blk00000001_sig00000519 : STD_LOGIC; 
  signal blk00000001_sig00000518 : STD_LOGIC; 
  signal blk00000001_sig00000517 : STD_LOGIC; 
  signal blk00000001_sig00000516 : STD_LOGIC; 
  signal blk00000001_sig00000515 : STD_LOGIC; 
  signal blk00000001_sig00000514 : STD_LOGIC; 
  signal blk00000001_sig00000513 : STD_LOGIC; 
  signal blk00000001_sig00000512 : STD_LOGIC; 
  signal blk00000001_sig00000511 : STD_LOGIC; 
  signal blk00000001_sig00000510 : STD_LOGIC; 
  signal blk00000001_sig0000050f : STD_LOGIC; 
  signal blk00000001_sig0000050e : STD_LOGIC; 
  signal blk00000001_sig0000050d : STD_LOGIC; 
  signal blk00000001_sig0000050c : STD_LOGIC; 
  signal blk00000001_sig0000050b : STD_LOGIC; 
  signal blk00000001_sig0000050a : STD_LOGIC; 
  signal blk00000001_sig00000509 : STD_LOGIC; 
  signal blk00000001_sig00000508 : STD_LOGIC; 
  signal blk00000001_sig00000507 : STD_LOGIC; 
  signal blk00000001_sig00000506 : STD_LOGIC; 
  signal blk00000001_sig00000505 : STD_LOGIC; 
  signal blk00000001_sig00000504 : STD_LOGIC; 
  signal blk00000001_sig00000503 : STD_LOGIC; 
  signal blk00000001_sig00000502 : STD_LOGIC; 
  signal blk00000001_sig00000501 : STD_LOGIC; 
  signal blk00000001_sig00000500 : STD_LOGIC; 
  signal blk00000001_sig000004ff : STD_LOGIC; 
  signal blk00000001_sig000004fe : STD_LOGIC; 
  signal blk00000001_sig000004fd : STD_LOGIC; 
  signal blk00000001_sig000004fc : STD_LOGIC; 
  signal blk00000001_sig000004fb : STD_LOGIC; 
  signal blk00000001_sig000004fa : STD_LOGIC; 
  signal blk00000001_sig000004f9 : STD_LOGIC; 
  signal blk00000001_sig000004f8 : STD_LOGIC; 
  signal blk00000001_sig000004f7 : STD_LOGIC; 
  signal blk00000001_sig000004f6 : STD_LOGIC; 
  signal blk00000001_sig000004f5 : STD_LOGIC; 
  signal blk00000001_sig000004f4 : STD_LOGIC; 
  signal blk00000001_sig000004f3 : STD_LOGIC; 
  signal blk00000001_sig000004f2 : STD_LOGIC; 
  signal blk00000001_sig000004f1 : STD_LOGIC; 
  signal blk00000001_sig000004f0 : STD_LOGIC; 
  signal blk00000001_sig000004ef : STD_LOGIC; 
  signal blk00000001_sig000004ee : STD_LOGIC; 
  signal blk00000001_sig000004ed : STD_LOGIC; 
  signal blk00000001_sig000004ec : STD_LOGIC; 
  signal blk00000001_sig000004eb : STD_LOGIC; 
  signal blk00000001_sig000004ea : STD_LOGIC; 
  signal blk00000001_sig000004e9 : STD_LOGIC; 
  signal blk00000001_sig000004e8 : STD_LOGIC; 
  signal blk00000001_sig000004e7 : STD_LOGIC; 
  signal blk00000001_sig000004e6 : STD_LOGIC; 
  signal blk00000001_sig000004e5 : STD_LOGIC; 
  signal blk00000001_sig000004e4 : STD_LOGIC; 
  signal blk00000001_sig000004e3 : STD_LOGIC; 
  signal blk00000001_sig000004e2 : STD_LOGIC; 
  signal blk00000001_sig000004e1 : STD_LOGIC; 
  signal blk00000001_sig000004e0 : STD_LOGIC; 
  signal blk00000001_sig000004df : STD_LOGIC; 
  signal blk00000001_sig000004de : STD_LOGIC; 
  signal blk00000001_sig000004dd : STD_LOGIC; 
  signal blk00000001_sig000004dc : STD_LOGIC; 
  signal blk00000001_sig000004db : STD_LOGIC; 
  signal blk00000001_sig000004da : STD_LOGIC; 
  signal blk00000001_sig000004d9 : STD_LOGIC; 
  signal blk00000001_sig000004d8 : STD_LOGIC; 
  signal blk00000001_sig000004d7 : STD_LOGIC; 
  signal blk00000001_sig000004d6 : STD_LOGIC; 
  signal blk00000001_sig000004d5 : STD_LOGIC; 
  signal blk00000001_sig000004d4 : STD_LOGIC; 
  signal blk00000001_sig000004d3 : STD_LOGIC; 
  signal blk00000001_sig000004d2 : STD_LOGIC; 
  signal blk00000001_sig000004d1 : STD_LOGIC; 
  signal blk00000001_sig000004d0 : STD_LOGIC; 
  signal blk00000001_sig000004cf : STD_LOGIC; 
  signal blk00000001_sig000004ce : STD_LOGIC; 
  signal blk00000001_sig000004cd : STD_LOGIC; 
  signal blk00000001_sig000004cc : STD_LOGIC; 
  signal blk00000001_sig000004cb : STD_LOGIC; 
  signal blk00000001_sig000004ca : STD_LOGIC; 
  signal blk00000001_sig000004c9 : STD_LOGIC; 
  signal blk00000001_sig000004c8 : STD_LOGIC; 
  signal blk00000001_sig000004c7 : STD_LOGIC; 
  signal blk00000001_sig000004c6 : STD_LOGIC; 
  signal blk00000001_sig000004c5 : STD_LOGIC; 
  signal blk00000001_sig000004c4 : STD_LOGIC; 
  signal blk00000001_sig000004c3 : STD_LOGIC; 
  signal blk00000001_sig000004c2 : STD_LOGIC; 
  signal blk00000001_sig000004c1 : STD_LOGIC; 
  signal blk00000001_sig000004c0 : STD_LOGIC; 
  signal blk00000001_sig000004bf : STD_LOGIC; 
  signal blk00000001_sig000004be : STD_LOGIC; 
  signal blk00000001_sig000004bd : STD_LOGIC; 
  signal blk00000001_sig000004bc : STD_LOGIC; 
  signal blk00000001_sig000004bb : STD_LOGIC; 
  signal blk00000001_sig000004ba : STD_LOGIC; 
  signal blk00000001_sig000004b9 : STD_LOGIC; 
  signal blk00000001_sig000004b8 : STD_LOGIC; 
  signal blk00000001_sig000004b7 : STD_LOGIC; 
  signal blk00000001_sig000004b6 : STD_LOGIC; 
  signal blk00000001_sig000004b5 : STD_LOGIC; 
  signal blk00000001_sig000004b4 : STD_LOGIC; 
  signal blk00000001_sig000004b3 : STD_LOGIC; 
  signal blk00000001_sig000004b2 : STD_LOGIC; 
  signal blk00000001_sig000004b1 : STD_LOGIC; 
  signal blk00000001_sig000004b0 : STD_LOGIC; 
  signal blk00000001_sig000004af : STD_LOGIC; 
  signal blk00000001_sig000004ae : STD_LOGIC; 
  signal blk00000001_sig000004ad : STD_LOGIC; 
  signal blk00000001_sig000004ac : STD_LOGIC; 
  signal blk00000001_sig000004ab : STD_LOGIC; 
  signal blk00000001_sig000004aa : STD_LOGIC; 
  signal blk00000001_sig000004a9 : STD_LOGIC; 
  signal blk00000001_sig000004a8 : STD_LOGIC; 
  signal blk00000001_sig000004a7 : STD_LOGIC; 
  signal blk00000001_sig000004a6 : STD_LOGIC; 
  signal blk00000001_sig000004a5 : STD_LOGIC; 
  signal blk00000001_sig000004a4 : STD_LOGIC; 
  signal blk00000001_sig000004a3 : STD_LOGIC; 
  signal blk00000001_sig000004a2 : STD_LOGIC; 
  signal blk00000001_sig000004a1 : STD_LOGIC; 
  signal blk00000001_sig000004a0 : STD_LOGIC; 
  signal blk00000001_sig0000049f : STD_LOGIC; 
  signal blk00000001_sig0000049e : STD_LOGIC; 
  signal blk00000001_sig0000049d : STD_LOGIC; 
  signal blk00000001_sig0000049c : STD_LOGIC; 
  signal blk00000001_sig0000049b : STD_LOGIC; 
  signal blk00000001_sig0000049a : STD_LOGIC; 
  signal blk00000001_sig00000499 : STD_LOGIC; 
  signal blk00000001_sig00000498 : STD_LOGIC; 
  signal blk00000001_sig00000497 : STD_LOGIC; 
  signal blk00000001_sig00000496 : STD_LOGIC; 
  signal blk00000001_sig00000495 : STD_LOGIC; 
  signal blk00000001_sig00000494 : STD_LOGIC; 
  signal blk00000001_sig00000493 : STD_LOGIC; 
  signal blk00000001_sig00000492 : STD_LOGIC; 
  signal blk00000001_sig00000491 : STD_LOGIC; 
  signal blk00000001_sig00000490 : STD_LOGIC; 
  signal blk00000001_sig0000048f : STD_LOGIC; 
  signal blk00000001_sig0000048e : STD_LOGIC; 
  signal blk00000001_sig0000048d : STD_LOGIC; 
  signal blk00000001_sig0000048c : STD_LOGIC; 
  signal blk00000001_sig0000048b : STD_LOGIC; 
  signal blk00000001_sig0000048a : STD_LOGIC; 
  signal blk00000001_sig00000489 : STD_LOGIC; 
  signal blk00000001_sig00000488 : STD_LOGIC; 
  signal blk00000001_sig00000487 : STD_LOGIC; 
  signal blk00000001_sig00000486 : STD_LOGIC; 
  signal blk00000001_sig00000485 : STD_LOGIC; 
  signal blk00000001_sig00000484 : STD_LOGIC; 
  signal blk00000001_sig00000483 : STD_LOGIC; 
  signal blk00000001_sig00000482 : STD_LOGIC; 
  signal blk00000001_sig00000481 : STD_LOGIC; 
  signal blk00000001_sig00000480 : STD_LOGIC; 
  signal blk00000001_sig0000047f : STD_LOGIC; 
  signal blk00000001_sig0000047e : STD_LOGIC; 
  signal blk00000001_sig0000047d : STD_LOGIC; 
  signal blk00000001_sig0000047c : STD_LOGIC; 
  signal blk00000001_sig0000047b : STD_LOGIC; 
  signal blk00000001_sig0000047a : STD_LOGIC; 
  signal blk00000001_sig00000479 : STD_LOGIC; 
  signal blk00000001_sig00000478 : STD_LOGIC; 
  signal blk00000001_sig00000477 : STD_LOGIC; 
  signal blk00000001_sig00000476 : STD_LOGIC; 
  signal blk00000001_sig00000475 : STD_LOGIC; 
  signal blk00000001_sig00000474 : STD_LOGIC; 
  signal blk00000001_sig00000473 : STD_LOGIC; 
  signal blk00000001_sig00000472 : STD_LOGIC; 
  signal blk00000001_sig00000471 : STD_LOGIC; 
  signal blk00000001_sig00000470 : STD_LOGIC; 
  signal blk00000001_sig0000046f : STD_LOGIC; 
  signal blk00000001_sig0000046e : STD_LOGIC; 
  signal blk00000001_sig0000046d : STD_LOGIC; 
  signal blk00000001_sig0000046c : STD_LOGIC; 
  signal blk00000001_sig0000046b : STD_LOGIC; 
  signal blk00000001_sig0000046a : STD_LOGIC; 
  signal blk00000001_sig00000469 : STD_LOGIC; 
  signal blk00000001_sig00000468 : STD_LOGIC; 
  signal blk00000001_sig00000467 : STD_LOGIC; 
  signal blk00000001_sig00000466 : STD_LOGIC; 
  signal blk00000001_sig00000465 : STD_LOGIC; 
  signal blk00000001_sig00000464 : STD_LOGIC; 
  signal blk00000001_sig00000463 : STD_LOGIC; 
  signal blk00000001_sig00000462 : STD_LOGIC; 
  signal blk00000001_sig00000461 : STD_LOGIC; 
  signal blk00000001_sig00000460 : STD_LOGIC; 
  signal blk00000001_sig0000045f : STD_LOGIC; 
  signal blk00000001_sig0000045e : STD_LOGIC; 
  signal blk00000001_sig0000045d : STD_LOGIC; 
  signal blk00000001_sig0000045c : STD_LOGIC; 
  signal blk00000001_sig0000045b : STD_LOGIC; 
  signal blk00000001_sig0000045a : STD_LOGIC; 
  signal blk00000001_sig00000459 : STD_LOGIC; 
  signal blk00000001_sig00000458 : STD_LOGIC; 
  signal blk00000001_sig00000457 : STD_LOGIC; 
  signal blk00000001_sig00000456 : STD_LOGIC; 
  signal blk00000001_sig00000455 : STD_LOGIC; 
  signal blk00000001_sig00000454 : STD_LOGIC; 
  signal blk00000001_sig00000453 : STD_LOGIC; 
  signal blk00000001_sig00000452 : STD_LOGIC; 
  signal blk00000001_sig00000451 : STD_LOGIC; 
  signal blk00000001_sig00000450 : STD_LOGIC; 
  signal blk00000001_sig0000044f : STD_LOGIC; 
  signal blk00000001_sig0000044e : STD_LOGIC; 
  signal blk00000001_sig0000044d : STD_LOGIC; 
  signal blk00000001_sig0000044c : STD_LOGIC; 
  signal blk00000001_sig0000044b : STD_LOGIC; 
  signal blk00000001_sig0000044a : STD_LOGIC; 
  signal blk00000001_sig00000449 : STD_LOGIC; 
  signal blk00000001_sig00000448 : STD_LOGIC; 
  signal blk00000001_sig00000447 : STD_LOGIC; 
  signal blk00000001_sig00000446 : STD_LOGIC; 
  signal blk00000001_sig00000445 : STD_LOGIC; 
  signal blk00000001_sig00000444 : STD_LOGIC; 
  signal blk00000001_sig00000443 : STD_LOGIC; 
  signal blk00000001_sig00000442 : STD_LOGIC; 
  signal blk00000001_sig00000441 : STD_LOGIC; 
  signal blk00000001_sig00000440 : STD_LOGIC; 
  signal blk00000001_sig0000043f : STD_LOGIC; 
  signal blk00000001_sig0000043e : STD_LOGIC; 
  signal blk00000001_sig0000043d : STD_LOGIC; 
  signal blk00000001_sig0000043c : STD_LOGIC; 
  signal blk00000001_sig0000043b : STD_LOGIC; 
  signal blk00000001_sig0000043a : STD_LOGIC; 
  signal blk00000001_sig00000439 : STD_LOGIC; 
  signal blk00000001_sig00000438 : STD_LOGIC; 
  signal blk00000001_sig00000437 : STD_LOGIC; 
  signal blk00000001_sig00000436 : STD_LOGIC; 
  signal blk00000001_sig00000435 : STD_LOGIC; 
  signal blk00000001_sig00000434 : STD_LOGIC; 
  signal blk00000001_sig00000433 : STD_LOGIC; 
  signal blk00000001_sig00000432 : STD_LOGIC; 
  signal blk00000001_sig00000431 : STD_LOGIC; 
  signal blk00000001_sig00000430 : STD_LOGIC; 
  signal blk00000001_sig0000042f : STD_LOGIC; 
  signal blk00000001_sig0000042e : STD_LOGIC; 
  signal blk00000001_sig0000042d : STD_LOGIC; 
  signal blk00000001_sig0000042c : STD_LOGIC; 
  signal blk00000001_sig0000042b : STD_LOGIC; 
  signal blk00000001_sig0000042a : STD_LOGIC; 
  signal blk00000001_sig00000429 : STD_LOGIC; 
  signal blk00000001_sig00000428 : STD_LOGIC; 
  signal blk00000001_sig00000427 : STD_LOGIC; 
  signal blk00000001_sig00000426 : STD_LOGIC; 
  signal blk00000001_sig00000425 : STD_LOGIC; 
  signal blk00000001_sig00000424 : STD_LOGIC; 
  signal blk00000001_sig00000423 : STD_LOGIC; 
  signal blk00000001_sig00000422 : STD_LOGIC; 
  signal blk00000001_sig00000421 : STD_LOGIC; 
  signal blk00000001_sig00000420 : STD_LOGIC; 
  signal blk00000001_sig0000041f : STD_LOGIC; 
  signal blk00000001_sig0000041e : STD_LOGIC; 
  signal blk00000001_sig0000041d : STD_LOGIC; 
  signal blk00000001_sig0000041c : STD_LOGIC; 
  signal blk00000001_sig0000041b : STD_LOGIC; 
  signal blk00000001_sig0000041a : STD_LOGIC; 
  signal blk00000001_sig00000419 : STD_LOGIC; 
  signal blk00000001_sig00000418 : STD_LOGIC; 
  signal blk00000001_sig00000417 : STD_LOGIC; 
  signal blk00000001_sig00000416 : STD_LOGIC; 
  signal blk00000001_sig00000415 : STD_LOGIC; 
  signal blk00000001_sig00000414 : STD_LOGIC; 
  signal blk00000001_sig00000413 : STD_LOGIC; 
  signal blk00000001_sig00000412 : STD_LOGIC; 
  signal blk00000001_sig00000411 : STD_LOGIC; 
  signal blk00000001_sig00000410 : STD_LOGIC; 
  signal blk00000001_sig0000040f : STD_LOGIC; 
  signal blk00000001_sig0000040e : STD_LOGIC; 
  signal blk00000001_sig0000040d : STD_LOGIC; 
  signal blk00000001_sig0000040c : STD_LOGIC; 
  signal blk00000001_sig0000040b : STD_LOGIC; 
  signal blk00000001_sig0000040a : STD_LOGIC; 
  signal blk00000001_sig00000409 : STD_LOGIC; 
  signal blk00000001_sig00000408 : STD_LOGIC; 
  signal blk00000001_sig00000407 : STD_LOGIC; 
  signal blk00000001_sig00000406 : STD_LOGIC; 
  signal blk00000001_sig00000405 : STD_LOGIC; 
  signal blk00000001_sig00000404 : STD_LOGIC; 
  signal blk00000001_sig00000403 : STD_LOGIC; 
  signal blk00000001_sig00000402 : STD_LOGIC; 
  signal blk00000001_sig00000401 : STD_LOGIC; 
  signal blk00000001_sig00000400 : STD_LOGIC; 
  signal blk00000001_sig000003ff : STD_LOGIC; 
  signal blk00000001_sig000003fe : STD_LOGIC; 
  signal blk00000001_sig000003fd : STD_LOGIC; 
  signal blk00000001_sig000003fc : STD_LOGIC; 
  signal blk00000001_sig000003fb : STD_LOGIC; 
  signal blk00000001_sig000003fa : STD_LOGIC; 
  signal blk00000001_sig000003f9 : STD_LOGIC; 
  signal blk00000001_sig000003f8 : STD_LOGIC; 
  signal blk00000001_sig000003f7 : STD_LOGIC; 
  signal blk00000001_sig000003f6 : STD_LOGIC; 
  signal blk00000001_sig000003f5 : STD_LOGIC; 
  signal blk00000001_sig000003f4 : STD_LOGIC; 
  signal blk00000001_sig000003f3 : STD_LOGIC; 
  signal blk00000001_sig000003f2 : STD_LOGIC; 
  signal blk00000001_sig000003f1 : STD_LOGIC; 
  signal blk00000001_sig000003f0 : STD_LOGIC; 
  signal blk00000001_sig000003ef : STD_LOGIC; 
  signal blk00000001_sig000003ee : STD_LOGIC; 
  signal blk00000001_sig000003ed : STD_LOGIC; 
  signal blk00000001_sig000003ec : STD_LOGIC; 
  signal blk00000001_sig000003eb : STD_LOGIC; 
  signal blk00000001_sig000003ea : STD_LOGIC; 
  signal blk00000001_sig000003e9 : STD_LOGIC; 
  signal blk00000001_sig000003e8 : STD_LOGIC; 
  signal blk00000001_sig000003e7 : STD_LOGIC; 
  signal blk00000001_sig000003e6 : STD_LOGIC; 
  signal blk00000001_sig000003e5 : STD_LOGIC; 
  signal blk00000001_sig000003e4 : STD_LOGIC; 
  signal blk00000001_sig000003e3 : STD_LOGIC; 
  signal blk00000001_sig000003e2 : STD_LOGIC; 
  signal blk00000001_sig000003e1 : STD_LOGIC; 
  signal blk00000001_sig000003e0 : STD_LOGIC; 
  signal blk00000001_sig000003df : STD_LOGIC; 
  signal blk00000001_sig000003de : STD_LOGIC; 
  signal blk00000001_sig000003dd : STD_LOGIC; 
  signal blk00000001_sig000003dc : STD_LOGIC; 
  signal blk00000001_sig000003db : STD_LOGIC; 
  signal blk00000001_sig000003da : STD_LOGIC; 
  signal blk00000001_sig000003d9 : STD_LOGIC; 
  signal blk00000001_sig000003d8 : STD_LOGIC; 
  signal blk00000001_sig000003d7 : STD_LOGIC; 
  signal blk00000001_sig000003d6 : STD_LOGIC; 
  signal blk00000001_sig000003d5 : STD_LOGIC; 
  signal blk00000001_sig000003d4 : STD_LOGIC; 
  signal blk00000001_sig000003d3 : STD_LOGIC; 
  signal blk00000001_sig000003d2 : STD_LOGIC; 
  signal blk00000001_sig000003d1 : STD_LOGIC; 
  signal blk00000001_sig000003d0 : STD_LOGIC; 
  signal blk00000001_sig000003cf : STD_LOGIC; 
  signal blk00000001_sig000003ce : STD_LOGIC; 
  signal blk00000001_sig000003cd : STD_LOGIC; 
  signal blk00000001_sig000003cc : STD_LOGIC; 
  signal blk00000001_sig000003cb : STD_LOGIC; 
  signal blk00000001_sig000003ca : STD_LOGIC; 
  signal blk00000001_sig000003c9 : STD_LOGIC; 
  signal blk00000001_sig000003c8 : STD_LOGIC; 
  signal blk00000001_sig000003c7 : STD_LOGIC; 
  signal blk00000001_sig000003c6 : STD_LOGIC; 
  signal blk00000001_sig000003c5 : STD_LOGIC; 
  signal blk00000001_sig000003c4 : STD_LOGIC; 
  signal blk00000001_sig000003c3 : STD_LOGIC; 
  signal blk00000001_sig000003c2 : STD_LOGIC; 
  signal blk00000001_sig000003c1 : STD_LOGIC; 
  signal blk00000001_sig000003c0 : STD_LOGIC; 
  signal blk00000001_sig000003bf : STD_LOGIC; 
  signal blk00000001_sig000003be : STD_LOGIC; 
  signal blk00000001_sig000003bd : STD_LOGIC; 
  signal blk00000001_sig000003bc : STD_LOGIC; 
  signal blk00000001_sig000003bb : STD_LOGIC; 
  signal blk00000001_sig000003ba : STD_LOGIC; 
  signal blk00000001_sig000003b9 : STD_LOGIC; 
  signal blk00000001_sig000003b8 : STD_LOGIC; 
  signal blk00000001_sig000003b7 : STD_LOGIC; 
  signal blk00000001_sig000003b6 : STD_LOGIC; 
  signal blk00000001_sig000003b5 : STD_LOGIC; 
  signal blk00000001_sig000003b4 : STD_LOGIC; 
  signal blk00000001_sig000003b3 : STD_LOGIC; 
  signal blk00000001_sig000003b2 : STD_LOGIC; 
  signal blk00000001_sig000003b1 : STD_LOGIC; 
  signal blk00000001_sig000003b0 : STD_LOGIC; 
  signal blk00000001_sig000003af : STD_LOGIC; 
  signal blk00000001_sig000003ae : STD_LOGIC; 
  signal blk00000001_sig000003ad : STD_LOGIC; 
  signal blk00000001_sig000003ac : STD_LOGIC; 
  signal blk00000001_sig000003ab : STD_LOGIC; 
  signal blk00000001_sig000003aa : STD_LOGIC; 
  signal blk00000001_sig000003a9 : STD_LOGIC; 
  signal blk00000001_sig000003a8 : STD_LOGIC; 
  signal blk00000001_sig000003a7 : STD_LOGIC; 
  signal blk00000001_sig000003a6 : STD_LOGIC; 
  signal blk00000001_sig000003a5 : STD_LOGIC; 
  signal blk00000001_sig000003a4 : STD_LOGIC; 
  signal blk00000001_sig000003a3 : STD_LOGIC; 
  signal blk00000001_sig000003a2 : STD_LOGIC; 
  signal blk00000001_sig000003a1 : STD_LOGIC; 
  signal blk00000001_sig000003a0 : STD_LOGIC; 
  signal blk00000001_sig0000039f : STD_LOGIC; 
  signal blk00000001_sig0000039e : STD_LOGIC; 
  signal blk00000001_sig0000039d : STD_LOGIC; 
  signal blk00000001_sig0000039c : STD_LOGIC; 
  signal blk00000001_sig0000039b : STD_LOGIC; 
  signal blk00000001_sig0000039a : STD_LOGIC; 
  signal blk00000001_sig00000399 : STD_LOGIC; 
  signal blk00000001_sig00000398 : STD_LOGIC; 
  signal blk00000001_sig00000397 : STD_LOGIC; 
  signal blk00000001_sig00000396 : STD_LOGIC; 
  signal blk00000001_sig00000395 : STD_LOGIC; 
  signal blk00000001_sig00000394 : STD_LOGIC; 
  signal blk00000001_sig00000393 : STD_LOGIC; 
  signal blk00000001_sig00000392 : STD_LOGIC; 
  signal blk00000001_sig00000391 : STD_LOGIC; 
  signal blk00000001_sig00000390 : STD_LOGIC; 
  signal blk00000001_sig0000038f : STD_LOGIC; 
  signal blk00000001_sig0000038e : STD_LOGIC; 
  signal blk00000001_sig0000038d : STD_LOGIC; 
  signal blk00000001_sig0000038c : STD_LOGIC; 
  signal blk00000001_sig0000038b : STD_LOGIC; 
  signal blk00000001_sig0000038a : STD_LOGIC; 
  signal blk00000001_sig00000389 : STD_LOGIC; 
  signal blk00000001_sig00000388 : STD_LOGIC; 
  signal blk00000001_sig00000387 : STD_LOGIC; 
  signal blk00000001_sig00000386 : STD_LOGIC; 
  signal blk00000001_sig00000385 : STD_LOGIC; 
  signal blk00000001_sig00000384 : STD_LOGIC; 
  signal blk00000001_sig00000383 : STD_LOGIC; 
  signal blk00000001_sig00000382 : STD_LOGIC; 
  signal blk00000001_sig00000381 : STD_LOGIC; 
  signal blk00000001_sig00000380 : STD_LOGIC; 
  signal blk00000001_sig0000037f : STD_LOGIC; 
  signal blk00000001_sig0000037e : STD_LOGIC; 
  signal blk00000001_sig0000037d : STD_LOGIC; 
  signal blk00000001_sig0000037c : STD_LOGIC; 
  signal blk00000001_sig0000037b : STD_LOGIC; 
  signal blk00000001_sig0000037a : STD_LOGIC; 
  signal blk00000001_sig00000379 : STD_LOGIC; 
  signal blk00000001_sig00000378 : STD_LOGIC; 
  signal blk00000001_sig00000377 : STD_LOGIC; 
  signal blk00000001_sig00000376 : STD_LOGIC; 
  signal blk00000001_sig00000375 : STD_LOGIC; 
  signal blk00000001_sig00000374 : STD_LOGIC; 
  signal blk00000001_sig00000373 : STD_LOGIC; 
  signal blk00000001_sig00000372 : STD_LOGIC; 
  signal blk00000001_sig00000371 : STD_LOGIC; 
  signal blk00000001_sig00000370 : STD_LOGIC; 
  signal blk00000001_sig0000036f : STD_LOGIC; 
  signal blk00000001_sig0000036e : STD_LOGIC; 
  signal blk00000001_sig0000036d : STD_LOGIC; 
  signal blk00000001_sig0000036c : STD_LOGIC; 
  signal blk00000001_sig0000036b : STD_LOGIC; 
  signal blk00000001_sig0000036a : STD_LOGIC; 
  signal blk00000001_sig00000369 : STD_LOGIC; 
  signal blk00000001_sig00000368 : STD_LOGIC; 
  signal blk00000001_sig00000367 : STD_LOGIC; 
  signal blk00000001_sig00000366 : STD_LOGIC; 
  signal blk00000001_sig00000365 : STD_LOGIC; 
  signal blk00000001_sig00000364 : STD_LOGIC; 
  signal blk00000001_sig00000363 : STD_LOGIC; 
  signal blk00000001_sig00000362 : STD_LOGIC; 
  signal blk00000001_sig00000361 : STD_LOGIC; 
  signal blk00000001_sig00000360 : STD_LOGIC; 
  signal blk00000001_sig0000035f : STD_LOGIC; 
  signal blk00000001_sig0000035e : STD_LOGIC; 
  signal blk00000001_sig0000035d : STD_LOGIC; 
  signal blk00000001_sig0000035c : STD_LOGIC; 
  signal blk00000001_sig0000035b : STD_LOGIC; 
  signal blk00000001_sig0000035a : STD_LOGIC; 
  signal blk00000001_sig00000359 : STD_LOGIC; 
  signal blk00000001_sig00000358 : STD_LOGIC; 
  signal blk00000001_sig00000357 : STD_LOGIC; 
  signal blk00000001_sig00000356 : STD_LOGIC; 
  signal blk00000001_sig00000355 : STD_LOGIC; 
  signal blk00000001_sig00000354 : STD_LOGIC; 
  signal blk00000001_sig00000353 : STD_LOGIC; 
  signal blk00000001_sig00000352 : STD_LOGIC; 
  signal blk00000001_sig00000351 : STD_LOGIC; 
  signal blk00000001_sig00000350 : STD_LOGIC; 
  signal blk00000001_sig0000034f : STD_LOGIC; 
  signal blk00000001_sig0000034e : STD_LOGIC; 
  signal blk00000001_sig0000034d : STD_LOGIC; 
  signal blk00000001_sig0000034c : STD_LOGIC; 
  signal blk00000001_sig0000034b : STD_LOGIC; 
  signal blk00000001_sig0000034a : STD_LOGIC; 
  signal blk00000001_sig00000349 : STD_LOGIC; 
  signal blk00000001_sig00000348 : STD_LOGIC; 
  signal blk00000001_sig00000347 : STD_LOGIC; 
  signal blk00000001_sig00000346 : STD_LOGIC; 
  signal blk00000001_sig00000345 : STD_LOGIC; 
  signal blk00000001_sig00000344 : STD_LOGIC; 
  signal blk00000001_sig00000343 : STD_LOGIC; 
  signal blk00000001_sig00000342 : STD_LOGIC; 
  signal blk00000001_sig00000341 : STD_LOGIC; 
  signal blk00000001_sig00000340 : STD_LOGIC; 
  signal blk00000001_sig0000033f : STD_LOGIC; 
  signal blk00000001_sig0000033e : STD_LOGIC; 
  signal blk00000001_sig0000033d : STD_LOGIC; 
  signal blk00000001_sig0000033c : STD_LOGIC; 
  signal blk00000001_sig0000033b : STD_LOGIC; 
  signal blk00000001_sig0000033a : STD_LOGIC; 
  signal blk00000001_sig00000339 : STD_LOGIC; 
  signal blk00000001_sig00000338 : STD_LOGIC; 
  signal blk00000001_sig00000337 : STD_LOGIC; 
  signal blk00000001_sig00000336 : STD_LOGIC; 
  signal blk00000001_sig00000335 : STD_LOGIC; 
  signal blk00000001_sig00000334 : STD_LOGIC; 
  signal blk00000001_sig00000333 : STD_LOGIC; 
  signal blk00000001_sig00000332 : STD_LOGIC; 
  signal blk00000001_sig00000331 : STD_LOGIC; 
  signal blk00000001_sig00000330 : STD_LOGIC; 
  signal blk00000001_sig0000032f : STD_LOGIC; 
  signal blk00000001_sig0000032e : STD_LOGIC; 
  signal blk00000001_sig0000032d : STD_LOGIC; 
  signal blk00000001_sig0000032c : STD_LOGIC; 
  signal blk00000001_sig0000032b : STD_LOGIC; 
  signal blk00000001_sig0000032a : STD_LOGIC; 
  signal blk00000001_sig00000329 : STD_LOGIC; 
  signal blk00000001_sig00000328 : STD_LOGIC; 
  signal blk00000001_sig00000327 : STD_LOGIC; 
  signal blk00000001_sig00000326 : STD_LOGIC; 
  signal blk00000001_sig00000325 : STD_LOGIC; 
  signal blk00000001_sig00000324 : STD_LOGIC; 
  signal blk00000001_sig00000323 : STD_LOGIC; 
  signal blk00000001_sig00000322 : STD_LOGIC; 
  signal blk00000001_sig00000321 : STD_LOGIC; 
  signal blk00000001_sig00000320 : STD_LOGIC; 
  signal blk00000001_sig0000031f : STD_LOGIC; 
  signal blk00000001_sig0000031e : STD_LOGIC; 
  signal blk00000001_sig0000031d : STD_LOGIC; 
  signal blk00000001_sig0000031c : STD_LOGIC; 
  signal blk00000001_sig0000031b : STD_LOGIC; 
  signal blk00000001_sig0000031a : STD_LOGIC; 
  signal blk00000001_sig00000319 : STD_LOGIC; 
  signal blk00000001_sig00000318 : STD_LOGIC; 
  signal blk00000001_sig00000317 : STD_LOGIC; 
  signal blk00000001_sig00000316 : STD_LOGIC; 
  signal blk00000001_sig00000315 : STD_LOGIC; 
  signal blk00000001_sig00000314 : STD_LOGIC; 
  signal blk00000001_sig00000313 : STD_LOGIC; 
  signal blk00000001_sig00000312 : STD_LOGIC; 
  signal blk00000001_sig00000311 : STD_LOGIC; 
  signal blk00000001_sig00000310 : STD_LOGIC; 
  signal blk00000001_sig0000030f : STD_LOGIC; 
  signal blk00000001_sig0000030e : STD_LOGIC; 
  signal blk00000001_sig0000030d : STD_LOGIC; 
  signal blk00000001_sig0000030c : STD_LOGIC; 
  signal blk00000001_sig0000030b : STD_LOGIC; 
  signal blk00000001_sig0000030a : STD_LOGIC; 
  signal blk00000001_sig00000309 : STD_LOGIC; 
  signal blk00000001_sig00000308 : STD_LOGIC; 
  signal blk00000001_sig00000307 : STD_LOGIC; 
  signal blk00000001_sig00000306 : STD_LOGIC; 
  signal blk00000001_sig00000305 : STD_LOGIC; 
  signal blk00000001_sig00000304 : STD_LOGIC; 
  signal blk00000001_sig00000303 : STD_LOGIC; 
  signal blk00000001_sig00000302 : STD_LOGIC; 
  signal blk00000001_sig00000301 : STD_LOGIC; 
  signal blk00000001_sig00000300 : STD_LOGIC; 
  signal blk00000001_sig000002ff : STD_LOGIC; 
  signal blk00000001_sig000002fe : STD_LOGIC; 
  signal blk00000001_sig000002fd : STD_LOGIC; 
  signal blk00000001_sig000002fc : STD_LOGIC; 
  signal blk00000001_sig000002fb : STD_LOGIC; 
  signal blk00000001_sig000002fa : STD_LOGIC; 
  signal blk00000001_sig000002f9 : STD_LOGIC; 
  signal blk00000001_sig000002f8 : STD_LOGIC; 
  signal blk00000001_sig000002f7 : STD_LOGIC; 
  signal blk00000001_sig000002f6 : STD_LOGIC; 
  signal blk00000001_sig000002f5 : STD_LOGIC; 
  signal blk00000001_sig000002f4 : STD_LOGIC; 
  signal blk00000001_sig000002f3 : STD_LOGIC; 
  signal blk00000001_sig000002f2 : STD_LOGIC; 
  signal blk00000001_sig000002f1 : STD_LOGIC; 
  signal blk00000001_sig000002f0 : STD_LOGIC; 
  signal blk00000001_sig000002ef : STD_LOGIC; 
  signal blk00000001_sig000002ee : STD_LOGIC; 
  signal blk00000001_sig000002ed : STD_LOGIC; 
  signal blk00000001_sig000002ec : STD_LOGIC; 
  signal blk00000001_sig000002eb : STD_LOGIC; 
  signal blk00000001_sig000002ea : STD_LOGIC; 
  signal blk00000001_sig000002e9 : STD_LOGIC; 
  signal blk00000001_sig000002e8 : STD_LOGIC; 
  signal blk00000001_sig000002e7 : STD_LOGIC; 
  signal blk00000001_sig000002e6 : STD_LOGIC; 
  signal blk00000001_sig000002e5 : STD_LOGIC; 
  signal blk00000001_sig000002e4 : STD_LOGIC; 
  signal blk00000001_sig000002e3 : STD_LOGIC; 
  signal blk00000001_sig000002e2 : STD_LOGIC; 
  signal blk00000001_sig000002e1 : STD_LOGIC; 
  signal blk00000001_sig000002e0 : STD_LOGIC; 
  signal blk00000001_sig000002df : STD_LOGIC; 
  signal blk00000001_sig000002de : STD_LOGIC; 
  signal blk00000001_sig000002dd : STD_LOGIC; 
  signal blk00000001_sig000002dc : STD_LOGIC; 
  signal blk00000001_sig000002db : STD_LOGIC; 
  signal blk00000001_sig000002da : STD_LOGIC; 
  signal blk00000001_sig000002d9 : STD_LOGIC; 
  signal blk00000001_sig000002d8 : STD_LOGIC; 
  signal blk00000001_sig000002d7 : STD_LOGIC; 
  signal blk00000001_sig000002d6 : STD_LOGIC; 
  signal blk00000001_sig000002d5 : STD_LOGIC; 
  signal blk00000001_sig000002d4 : STD_LOGIC; 
  signal blk00000001_sig000002d3 : STD_LOGIC; 
  signal blk00000001_sig000002d2 : STD_LOGIC; 
  signal blk00000001_sig000002d1 : STD_LOGIC; 
  signal blk00000001_sig000002d0 : STD_LOGIC; 
  signal blk00000001_sig000002cf : STD_LOGIC; 
  signal blk00000001_sig000002ce : STD_LOGIC; 
  signal blk00000001_sig000002cd : STD_LOGIC; 
  signal blk00000001_sig000002cc : STD_LOGIC; 
  signal blk00000001_sig000002cb : STD_LOGIC; 
  signal blk00000001_sig000002ca : STD_LOGIC; 
  signal blk00000001_sig000002c9 : STD_LOGIC; 
  signal blk00000001_sig000002c8 : STD_LOGIC; 
  signal blk00000001_sig000002c7 : STD_LOGIC; 
  signal blk00000001_sig000002c6 : STD_LOGIC; 
  signal blk00000001_sig000002c5 : STD_LOGIC; 
  signal blk00000001_sig000002c4 : STD_LOGIC; 
  signal blk00000001_sig000002c3 : STD_LOGIC; 
  signal blk00000001_sig000002c2 : STD_LOGIC; 
  signal blk00000001_sig000002c1 : STD_LOGIC; 
  signal blk00000001_sig000002c0 : STD_LOGIC; 
  signal blk00000001_sig000002bf : STD_LOGIC; 
  signal blk00000001_sig000002be : STD_LOGIC; 
  signal blk00000001_sig000002bd : STD_LOGIC; 
  signal blk00000001_sig000002bc : STD_LOGIC; 
  signal blk00000001_sig000002bb : STD_LOGIC; 
  signal blk00000001_sig000002ba : STD_LOGIC; 
  signal blk00000001_sig000002b9 : STD_LOGIC; 
  signal blk00000001_sig000002b8 : STD_LOGIC; 
  signal blk00000001_sig000002b7 : STD_LOGIC; 
  signal blk00000001_sig000002b6 : STD_LOGIC; 
  signal blk00000001_sig000002b5 : STD_LOGIC; 
  signal blk00000001_sig000002b4 : STD_LOGIC; 
  signal blk00000001_sig000002b3 : STD_LOGIC; 
  signal blk00000001_sig000002b2 : STD_LOGIC; 
  signal blk00000001_sig000002b1 : STD_LOGIC; 
  signal blk00000001_sig000002b0 : STD_LOGIC; 
  signal blk00000001_sig000002af : STD_LOGIC; 
  signal blk00000001_sig000002ae : STD_LOGIC; 
  signal blk00000001_sig000002ad : STD_LOGIC; 
  signal blk00000001_sig000002ac : STD_LOGIC; 
  signal blk00000001_sig000002ab : STD_LOGIC; 
  signal blk00000001_sig000002aa : STD_LOGIC; 
  signal blk00000001_sig000002a9 : STD_LOGIC; 
  signal blk00000001_sig000002a8 : STD_LOGIC; 
  signal blk00000001_sig000002a7 : STD_LOGIC; 
  signal blk00000001_sig000002a6 : STD_LOGIC; 
  signal blk00000001_sig000002a5 : STD_LOGIC; 
  signal blk00000001_sig000002a4 : STD_LOGIC; 
  signal blk00000001_sig000002a3 : STD_LOGIC; 
  signal blk00000001_sig000002a2 : STD_LOGIC; 
  signal blk00000001_sig000002a1 : STD_LOGIC; 
  signal blk00000001_sig000002a0 : STD_LOGIC; 
  signal blk00000001_sig0000029f : STD_LOGIC; 
  signal blk00000001_sig0000029e : STD_LOGIC; 
  signal blk00000001_sig0000029d : STD_LOGIC; 
  signal blk00000001_sig0000029c : STD_LOGIC; 
  signal blk00000001_sig0000029b : STD_LOGIC; 
  signal blk00000001_sig0000029a : STD_LOGIC; 
  signal blk00000001_sig00000299 : STD_LOGIC; 
  signal blk00000001_sig00000298 : STD_LOGIC; 
  signal blk00000001_sig00000297 : STD_LOGIC; 
  signal blk00000001_sig00000296 : STD_LOGIC; 
  signal blk00000001_sig00000295 : STD_LOGIC; 
  signal blk00000001_sig00000294 : STD_LOGIC; 
  signal blk00000001_sig00000293 : STD_LOGIC; 
  signal blk00000001_sig00000292 : STD_LOGIC; 
  signal blk00000001_sig00000291 : STD_LOGIC; 
  signal blk00000001_sig00000290 : STD_LOGIC; 
  signal blk00000001_sig0000028f : STD_LOGIC; 
  signal blk00000001_sig0000028e : STD_LOGIC; 
  signal blk00000001_sig0000028d : STD_LOGIC; 
  signal blk00000001_sig0000028c : STD_LOGIC; 
  signal blk00000001_sig0000028b : STD_LOGIC; 
  signal blk00000001_sig0000028a : STD_LOGIC; 
  signal blk00000001_sig00000289 : STD_LOGIC; 
  signal blk00000001_sig00000288 : STD_LOGIC; 
  signal blk00000001_sig00000287 : STD_LOGIC; 
  signal blk00000001_sig00000286 : STD_LOGIC; 
  signal blk00000001_sig00000285 : STD_LOGIC; 
  signal blk00000001_sig00000284 : STD_LOGIC; 
  signal blk00000001_sig00000283 : STD_LOGIC; 
  signal blk00000001_sig00000282 : STD_LOGIC; 
  signal blk00000001_sig00000281 : STD_LOGIC; 
  signal blk00000001_sig00000280 : STD_LOGIC; 
  signal blk00000001_sig0000027f : STD_LOGIC; 
  signal blk00000001_sig0000027e : STD_LOGIC; 
  signal blk00000001_sig0000027d : STD_LOGIC; 
  signal blk00000001_sig0000027c : STD_LOGIC; 
  signal blk00000001_sig0000027b : STD_LOGIC; 
  signal blk00000001_sig0000027a : STD_LOGIC; 
  signal blk00000001_sig00000279 : STD_LOGIC; 
  signal blk00000001_sig00000278 : STD_LOGIC; 
  signal blk00000001_sig00000277 : STD_LOGIC; 
  signal blk00000001_sig00000276 : STD_LOGIC; 
  signal blk00000001_sig00000275 : STD_LOGIC; 
  signal blk00000001_sig00000274 : STD_LOGIC; 
  signal blk00000001_sig00000273 : STD_LOGIC; 
  signal blk00000001_sig00000272 : STD_LOGIC; 
  signal blk00000001_sig00000271 : STD_LOGIC; 
  signal blk00000001_sig00000270 : STD_LOGIC; 
  signal blk00000001_sig0000026f : STD_LOGIC; 
  signal blk00000001_sig0000026e : STD_LOGIC; 
  signal blk00000001_sig0000026d : STD_LOGIC; 
  signal blk00000001_sig0000026c : STD_LOGIC; 
  signal blk00000001_sig0000026b : STD_LOGIC; 
  signal blk00000001_sig0000026a : STD_LOGIC; 
  signal blk00000001_sig00000269 : STD_LOGIC; 
  signal blk00000001_sig00000268 : STD_LOGIC; 
  signal blk00000001_sig00000267 : STD_LOGIC; 
  signal blk00000001_sig00000266 : STD_LOGIC; 
  signal blk00000001_sig00000265 : STD_LOGIC; 
  signal blk00000001_sig00000264 : STD_LOGIC; 
  signal blk00000001_sig00000263 : STD_LOGIC; 
  signal blk00000001_sig00000262 : STD_LOGIC; 
  signal blk00000001_sig00000261 : STD_LOGIC; 
  signal blk00000001_sig00000260 : STD_LOGIC; 
  signal blk00000001_sig0000025f : STD_LOGIC; 
  signal blk00000001_sig0000025e : STD_LOGIC; 
  signal blk00000001_sig0000025d : STD_LOGIC; 
  signal blk00000001_sig0000025c : STD_LOGIC; 
  signal blk00000001_sig0000025b : STD_LOGIC; 
  signal blk00000001_sig0000025a : STD_LOGIC; 
  signal blk00000001_sig00000259 : STD_LOGIC; 
  signal blk00000001_sig00000258 : STD_LOGIC; 
  signal blk00000001_sig00000257 : STD_LOGIC; 
  signal blk00000001_sig00000256 : STD_LOGIC; 
  signal blk00000001_sig00000255 : STD_LOGIC; 
  signal blk00000001_sig00000254 : STD_LOGIC; 
  signal blk00000001_sig00000253 : STD_LOGIC; 
  signal blk00000001_sig00000252 : STD_LOGIC; 
  signal blk00000001_sig00000251 : STD_LOGIC; 
  signal blk00000001_sig00000250 : STD_LOGIC; 
  signal blk00000001_sig0000024f : STD_LOGIC; 
  signal blk00000001_sig0000024e : STD_LOGIC; 
  signal blk00000001_sig0000024d : STD_LOGIC; 
  signal blk00000001_sig0000024c : STD_LOGIC; 
  signal blk00000001_sig0000024b : STD_LOGIC; 
  signal blk00000001_sig0000024a : STD_LOGIC; 
  signal blk00000001_sig00000249 : STD_LOGIC; 
  signal blk00000001_sig00000248 : STD_LOGIC; 
  signal blk00000001_sig00000247 : STD_LOGIC; 
  signal blk00000001_sig00000246 : STD_LOGIC; 
  signal blk00000001_sig00000245 : STD_LOGIC; 
  signal blk00000001_sig00000244 : STD_LOGIC; 
  signal blk00000001_sig00000243 : STD_LOGIC; 
  signal blk00000001_sig00000242 : STD_LOGIC; 
  signal blk00000001_sig00000241 : STD_LOGIC; 
  signal blk00000001_sig00000240 : STD_LOGIC; 
  signal blk00000001_sig0000023f : STD_LOGIC; 
  signal blk00000001_sig0000023e : STD_LOGIC; 
  signal blk00000001_sig0000023d : STD_LOGIC; 
  signal blk00000001_sig0000023c : STD_LOGIC; 
  signal blk00000001_sig0000023b : STD_LOGIC; 
  signal blk00000001_sig0000023a : STD_LOGIC; 
  signal blk00000001_sig00000239 : STD_LOGIC; 
  signal blk00000001_sig00000238 : STD_LOGIC; 
  signal blk00000001_sig00000237 : STD_LOGIC; 
  signal blk00000001_sig00000236 : STD_LOGIC; 
  signal blk00000001_sig00000235 : STD_LOGIC; 
  signal blk00000001_sig00000234 : STD_LOGIC; 
  signal blk00000001_sig00000233 : STD_LOGIC; 
  signal blk00000001_sig00000232 : STD_LOGIC; 
  signal blk00000001_sig00000231 : STD_LOGIC; 
  signal blk00000001_sig00000230 : STD_LOGIC; 
  signal blk00000001_sig0000022f : STD_LOGIC; 
  signal blk00000001_sig0000022e : STD_LOGIC; 
  signal blk00000001_sig0000022d : STD_LOGIC; 
  signal blk00000001_sig0000022c : STD_LOGIC; 
  signal blk00000001_sig0000022b : STD_LOGIC; 
  signal blk00000001_sig0000022a : STD_LOGIC; 
  signal blk00000001_sig00000229 : STD_LOGIC; 
  signal blk00000001_sig00000228 : STD_LOGIC; 
  signal blk00000001_sig00000227 : STD_LOGIC; 
  signal blk00000001_sig00000226 : STD_LOGIC; 
  signal blk00000001_sig00000225 : STD_LOGIC; 
  signal blk00000001_sig00000224 : STD_LOGIC; 
  signal blk00000001_sig00000223 : STD_LOGIC; 
  signal blk00000001_sig00000222 : STD_LOGIC; 
  signal blk00000001_sig00000221 : STD_LOGIC; 
  signal blk00000001_sig00000220 : STD_LOGIC; 
  signal blk00000001_sig0000021f : STD_LOGIC; 
  signal blk00000001_sig0000021e : STD_LOGIC; 
  signal blk00000001_sig0000021d : STD_LOGIC; 
  signal blk00000001_sig0000021c : STD_LOGIC; 
  signal blk00000001_sig0000021b : STD_LOGIC; 
  signal blk00000001_sig0000021a : STD_LOGIC; 
  signal blk00000001_sig00000219 : STD_LOGIC; 
  signal blk00000001_sig00000218 : STD_LOGIC; 
  signal blk00000001_sig00000217 : STD_LOGIC; 
  signal blk00000001_sig00000216 : STD_LOGIC; 
  signal blk00000001_sig00000215 : STD_LOGIC; 
  signal blk00000001_sig00000214 : STD_LOGIC; 
  signal blk00000001_sig00000213 : STD_LOGIC; 
  signal blk00000001_sig00000212 : STD_LOGIC; 
  signal blk00000001_sig00000211 : STD_LOGIC; 
  signal blk00000001_sig00000210 : STD_LOGIC; 
  signal blk00000001_sig0000020f : STD_LOGIC; 
  signal blk00000001_sig0000020e : STD_LOGIC; 
  signal blk00000001_sig0000020d : STD_LOGIC; 
  signal blk00000001_sig0000020c : STD_LOGIC; 
  signal blk00000001_sig0000020b : STD_LOGIC; 
  signal blk00000001_sig0000020a : STD_LOGIC; 
  signal blk00000001_sig00000209 : STD_LOGIC; 
  signal blk00000001_sig00000208 : STD_LOGIC; 
  signal blk00000001_sig00000207 : STD_LOGIC; 
  signal blk00000001_sig00000206 : STD_LOGIC; 
  signal blk00000001_sig00000205 : STD_LOGIC; 
  signal blk00000001_sig00000204 : STD_LOGIC; 
  signal blk00000001_sig00000203 : STD_LOGIC; 
  signal blk00000001_sig00000202 : STD_LOGIC; 
  signal blk00000001_sig00000201 : STD_LOGIC; 
  signal blk00000001_sig00000200 : STD_LOGIC; 
  signal blk00000001_sig000001ff : STD_LOGIC; 
  signal blk00000001_sig000001fe : STD_LOGIC; 
  signal blk00000001_sig000001fd : STD_LOGIC; 
  signal blk00000001_sig000001fc : STD_LOGIC; 
  signal blk00000001_sig000001fb : STD_LOGIC; 
  signal blk00000001_sig000001fa : STD_LOGIC; 
  signal blk00000001_sig000001f9 : STD_LOGIC; 
  signal blk00000001_sig000001f8 : STD_LOGIC; 
  signal blk00000001_sig000001f7 : STD_LOGIC; 
  signal blk00000001_sig000001f6 : STD_LOGIC; 
  signal blk00000001_sig000001f5 : STD_LOGIC; 
  signal blk00000001_sig000001f4 : STD_LOGIC; 
  signal blk00000001_sig000001f3 : STD_LOGIC; 
  signal blk00000001_sig000001f2 : STD_LOGIC; 
  signal blk00000001_sig000001f1 : STD_LOGIC; 
  signal blk00000001_sig000001f0 : STD_LOGIC; 
  signal blk00000001_sig000001ef : STD_LOGIC; 
  signal blk00000001_sig000001ee : STD_LOGIC; 
  signal blk00000001_sig000001ed : STD_LOGIC; 
  signal blk00000001_sig000001ec : STD_LOGIC; 
  signal blk00000001_sig000001eb : STD_LOGIC; 
  signal blk00000001_sig000001ea : STD_LOGIC; 
  signal blk00000001_sig000001e9 : STD_LOGIC; 
  signal blk00000001_sig000001e8 : STD_LOGIC; 
  signal blk00000001_sig000001e7 : STD_LOGIC; 
  signal blk00000001_sig000001e6 : STD_LOGIC; 
  signal blk00000001_sig000001e5 : STD_LOGIC; 
  signal blk00000001_sig000001e4 : STD_LOGIC; 
  signal blk00000001_sig000001e3 : STD_LOGIC; 
  signal blk00000001_sig000001e2 : STD_LOGIC; 
  signal blk00000001_sig000001e1 : STD_LOGIC; 
  signal blk00000001_sig000001e0 : STD_LOGIC; 
  signal blk00000001_sig000001df : STD_LOGIC; 
  signal blk00000001_sig000001de : STD_LOGIC; 
  signal blk00000001_sig000001dd : STD_LOGIC; 
  signal blk00000001_sig000001dc : STD_LOGIC; 
  signal blk00000001_sig000001db : STD_LOGIC; 
  signal blk00000001_sig000001da : STD_LOGIC; 
  signal blk00000001_sig000001d9 : STD_LOGIC; 
  signal blk00000001_sig000001d8 : STD_LOGIC; 
  signal blk00000001_sig000001d7 : STD_LOGIC; 
  signal blk00000001_sig000001d6 : STD_LOGIC; 
  signal blk00000001_sig000001d5 : STD_LOGIC; 
  signal blk00000001_sig000001d4 : STD_LOGIC; 
  signal blk00000001_sig000001d3 : STD_LOGIC; 
  signal blk00000001_sig000001d2 : STD_LOGIC; 
  signal blk00000001_sig000001d1 : STD_LOGIC; 
  signal blk00000001_sig000001d0 : STD_LOGIC; 
  signal blk00000001_sig000001cf : STD_LOGIC; 
  signal blk00000001_sig000001ce : STD_LOGIC; 
  signal blk00000001_sig000001cd : STD_LOGIC; 
  signal blk00000001_sig000001cc : STD_LOGIC; 
  signal blk00000001_sig000001cb : STD_LOGIC; 
  signal blk00000001_sig000001ca : STD_LOGIC; 
  signal blk00000001_sig000001c9 : STD_LOGIC; 
  signal blk00000001_sig000001c8 : STD_LOGIC; 
  signal blk00000001_sig000001c7 : STD_LOGIC; 
  signal blk00000001_sig000001c6 : STD_LOGIC; 
  signal blk00000001_sig000001c5 : STD_LOGIC; 
  signal blk00000001_sig000001c4 : STD_LOGIC; 
  signal blk00000001_sig000001c3 : STD_LOGIC; 
  signal blk00000001_sig000001c2 : STD_LOGIC; 
  signal blk00000001_sig000001c1 : STD_LOGIC; 
  signal blk00000001_sig000001c0 : STD_LOGIC; 
  signal blk00000001_sig000001bf : STD_LOGIC; 
  signal blk00000001_sig000001be : STD_LOGIC; 
  signal blk00000001_sig000001bd : STD_LOGIC; 
  signal blk00000001_sig000001bc : STD_LOGIC; 
  signal blk00000001_sig000001bb : STD_LOGIC; 
  signal blk00000001_sig000001ba : STD_LOGIC; 
  signal blk00000001_sig000001b9 : STD_LOGIC; 
  signal blk00000001_sig000001b8 : STD_LOGIC; 
  signal blk00000001_sig000001b7 : STD_LOGIC; 
  signal blk00000001_sig000001b6 : STD_LOGIC; 
  signal blk00000001_sig000001b5 : STD_LOGIC; 
  signal blk00000001_sig000001b4 : STD_LOGIC; 
  signal blk00000001_sig000001b3 : STD_LOGIC; 
  signal blk00000001_sig000001b2 : STD_LOGIC; 
  signal blk00000001_sig000001b1 : STD_LOGIC; 
  signal blk00000001_sig000001b0 : STD_LOGIC; 
  signal blk00000001_sig000001af : STD_LOGIC; 
  signal blk00000001_sig000001ae : STD_LOGIC; 
  signal blk00000001_sig000001ad : STD_LOGIC; 
  signal blk00000001_sig000001ac : STD_LOGIC; 
  signal blk00000001_sig000001ab : STD_LOGIC; 
  signal blk00000001_sig000001aa : STD_LOGIC; 
  signal blk00000001_sig000001a9 : STD_LOGIC; 
  signal blk00000001_sig000001a8 : STD_LOGIC; 
  signal blk00000001_sig000001a7 : STD_LOGIC; 
  signal blk00000001_sig000001a6 : STD_LOGIC; 
  signal blk00000001_sig000001a5 : STD_LOGIC; 
  signal blk00000001_sig000001a4 : STD_LOGIC; 
  signal blk00000001_sig000001a3 : STD_LOGIC; 
  signal blk00000001_sig000001a2 : STD_LOGIC; 
  signal blk00000001_sig000001a1 : STD_LOGIC; 
  signal blk00000001_sig000001a0 : STD_LOGIC; 
  signal blk00000001_sig0000019f : STD_LOGIC; 
  signal blk00000001_sig0000019e : STD_LOGIC; 
  signal blk00000001_sig0000019d : STD_LOGIC; 
  signal blk00000001_sig0000019c : STD_LOGIC; 
  signal blk00000001_sig0000019b : STD_LOGIC; 
  signal blk00000001_sig0000019a : STD_LOGIC; 
  signal blk00000001_sig00000199 : STD_LOGIC; 
  signal blk00000001_sig00000198 : STD_LOGIC; 
  signal blk00000001_sig00000197 : STD_LOGIC; 
  signal blk00000001_sig00000196 : STD_LOGIC; 
  signal blk00000001_sig00000195 : STD_LOGIC; 
  signal blk00000001_sig00000194 : STD_LOGIC; 
  signal blk00000001_sig00000193 : STD_LOGIC; 
  signal blk00000001_sig00000192 : STD_LOGIC; 
  signal blk00000001_sig00000191 : STD_LOGIC; 
  signal blk00000001_sig00000190 : STD_LOGIC; 
  signal blk00000001_sig0000018f : STD_LOGIC; 
  signal blk00000001_sig0000018e : STD_LOGIC; 
  signal blk00000001_sig0000018d : STD_LOGIC; 
  signal blk00000001_sig0000018c : STD_LOGIC; 
  signal blk00000001_sig0000018b : STD_LOGIC; 
  signal blk00000001_sig0000018a : STD_LOGIC; 
  signal blk00000001_sig00000189 : STD_LOGIC; 
  signal blk00000001_sig00000188 : STD_LOGIC; 
  signal blk00000001_sig00000187 : STD_LOGIC; 
  signal blk00000001_sig00000186 : STD_LOGIC; 
  signal blk00000001_sig00000185 : STD_LOGIC; 
  signal blk00000001_sig00000184 : STD_LOGIC; 
  signal blk00000001_sig00000183 : STD_LOGIC; 
  signal blk00000001_sig00000182 : STD_LOGIC; 
  signal blk00000001_sig00000181 : STD_LOGIC; 
  signal blk00000001_sig00000180 : STD_LOGIC; 
  signal blk00000001_sig0000017f : STD_LOGIC; 
  signal blk00000001_sig0000017e : STD_LOGIC; 
  signal blk00000001_sig0000017d : STD_LOGIC; 
  signal blk00000001_sig0000017c : STD_LOGIC; 
  signal blk00000001_sig0000017b : STD_LOGIC; 
  signal blk00000001_sig0000017a : STD_LOGIC; 
  signal blk00000001_sig00000179 : STD_LOGIC; 
  signal blk00000001_sig00000178 : STD_LOGIC; 
  signal blk00000001_sig00000177 : STD_LOGIC; 
  signal blk00000001_sig00000176 : STD_LOGIC; 
  signal blk00000001_sig00000175 : STD_LOGIC; 
  signal blk00000001_sig00000174 : STD_LOGIC; 
  signal blk00000001_sig00000173 : STD_LOGIC; 
  signal blk00000001_sig00000172 : STD_LOGIC; 
  signal blk00000001_sig00000171 : STD_LOGIC; 
  signal blk00000001_sig00000170 : STD_LOGIC; 
  signal blk00000001_sig0000016f : STD_LOGIC; 
  signal blk00000001_sig0000016e : STD_LOGIC; 
  signal blk00000001_sig0000016d : STD_LOGIC; 
  signal blk00000001_sig0000016c : STD_LOGIC; 
  signal blk00000001_sig0000016b : STD_LOGIC; 
  signal blk00000001_sig0000016a : STD_LOGIC; 
  signal blk00000001_sig00000169 : STD_LOGIC; 
  signal blk00000001_sig00000168 : STD_LOGIC; 
  signal blk00000001_sig00000167 : STD_LOGIC; 
  signal blk00000001_sig00000166 : STD_LOGIC; 
  signal blk00000001_sig00000165 : STD_LOGIC; 
  signal blk00000001_sig00000164 : STD_LOGIC; 
  signal blk00000001_sig00000163 : STD_LOGIC; 
  signal blk00000001_sig00000162 : STD_LOGIC; 
  signal blk00000001_sig00000161 : STD_LOGIC; 
  signal blk00000001_sig00000160 : STD_LOGIC; 
  signal blk00000001_sig0000015f : STD_LOGIC; 
  signal blk00000001_sig0000015e : STD_LOGIC; 
  signal blk00000001_sig0000015d : STD_LOGIC; 
  signal blk00000001_sig0000015c : STD_LOGIC; 
  signal blk00000001_sig0000015b : STD_LOGIC; 
  signal blk00000001_sig0000015a : STD_LOGIC; 
  signal blk00000001_sig00000159 : STD_LOGIC; 
  signal blk00000001_sig00000158 : STD_LOGIC; 
  signal blk00000001_sig00000157 : STD_LOGIC; 
  signal blk00000001_sig00000156 : STD_LOGIC; 
  signal blk00000001_sig00000155 : STD_LOGIC; 
  signal blk00000001_sig00000154 : STD_LOGIC; 
  signal blk00000001_sig00000153 : STD_LOGIC; 
  signal blk00000001_sig00000152 : STD_LOGIC; 
  signal blk00000001_sig00000151 : STD_LOGIC; 
  signal blk00000001_sig00000150 : STD_LOGIC; 
  signal blk00000001_sig0000014f : STD_LOGIC; 
  signal blk00000001_sig0000014e : STD_LOGIC; 
  signal blk00000001_sig0000014d : STD_LOGIC; 
  signal blk00000001_sig0000014c : STD_LOGIC; 
  signal blk00000001_sig0000014b : STD_LOGIC; 
  signal blk00000001_sig0000014a : STD_LOGIC; 
  signal blk00000001_sig00000149 : STD_LOGIC; 
  signal blk00000001_sig00000148 : STD_LOGIC; 
  signal blk00000001_sig00000147 : STD_LOGIC; 
  signal blk00000001_sig00000146 : STD_LOGIC; 
  signal blk00000001_sig00000145 : STD_LOGIC; 
  signal blk00000001_sig00000144 : STD_LOGIC; 
  signal blk00000001_sig00000143 : STD_LOGIC; 
  signal blk00000001_sig00000142 : STD_LOGIC; 
  signal blk00000001_sig00000141 : STD_LOGIC; 
  signal blk00000001_sig00000140 : STD_LOGIC; 
  signal blk00000001_sig0000013f : STD_LOGIC; 
  signal blk00000001_sig0000013e : STD_LOGIC; 
  signal blk00000001_sig0000013d : STD_LOGIC; 
  signal blk00000001_sig0000013c : STD_LOGIC; 
  signal blk00000001_sig0000013b : STD_LOGIC; 
  signal blk00000001_sig0000013a : STD_LOGIC; 
  signal blk00000001_sig00000139 : STD_LOGIC; 
  signal blk00000001_sig00000138 : STD_LOGIC; 
  signal blk00000001_sig00000137 : STD_LOGIC; 
  signal blk00000001_sig00000136 : STD_LOGIC; 
  signal blk00000001_sig00000135 : STD_LOGIC; 
  signal blk00000001_sig00000134 : STD_LOGIC; 
  signal blk00000001_sig00000133 : STD_LOGIC; 
  signal blk00000001_sig00000132 : STD_LOGIC; 
  signal blk00000001_sig00000131 : STD_LOGIC; 
  signal blk00000001_sig00000130 : STD_LOGIC; 
  signal blk00000001_sig0000012f : STD_LOGIC; 
  signal blk00000001_sig0000012e : STD_LOGIC; 
  signal blk00000001_sig0000012d : STD_LOGIC; 
  signal blk00000001_sig0000012c : STD_LOGIC; 
  signal blk00000001_sig0000012b : STD_LOGIC; 
  signal blk00000001_sig0000012a : STD_LOGIC; 
  signal blk00000001_sig00000129 : STD_LOGIC; 
  signal blk00000001_sig00000128 : STD_LOGIC; 
  signal blk00000001_sig00000127 : STD_LOGIC; 
  signal blk00000001_sig00000126 : STD_LOGIC; 
  signal blk00000001_sig00000125 : STD_LOGIC; 
  signal blk00000001_sig00000124 : STD_LOGIC; 
  signal blk00000001_sig00000123 : STD_LOGIC; 
  signal blk00000001_sig00000122 : STD_LOGIC; 
  signal blk00000001_sig00000121 : STD_LOGIC; 
  signal blk00000001_sig00000120 : STD_LOGIC; 
  signal blk00000001_sig0000011f : STD_LOGIC; 
  signal blk00000001_sig0000011e : STD_LOGIC; 
  signal blk00000001_sig0000011d : STD_LOGIC; 
  signal blk00000001_sig0000011c : STD_LOGIC; 
  signal blk00000001_sig0000011b : STD_LOGIC; 
  signal blk00000001_sig0000011a : STD_LOGIC; 
  signal blk00000001_sig00000119 : STD_LOGIC; 
  signal blk00000001_sig00000118 : STD_LOGIC; 
  signal blk00000001_sig00000117 : STD_LOGIC; 
  signal blk00000001_sig00000116 : STD_LOGIC; 
  signal blk00000001_sig00000115 : STD_LOGIC; 
  signal blk00000001_sig00000114 : STD_LOGIC; 
  signal blk00000001_sig00000113 : STD_LOGIC; 
  signal blk00000001_sig00000112 : STD_LOGIC; 
  signal blk00000001_sig00000111 : STD_LOGIC; 
  signal blk00000001_sig00000110 : STD_LOGIC; 
  signal blk00000001_sig0000010f : STD_LOGIC; 
  signal blk00000001_sig0000010e : STD_LOGIC; 
  signal blk00000001_sig0000010d : STD_LOGIC; 
  signal blk00000001_sig0000010c : STD_LOGIC; 
  signal blk00000001_sig0000010b : STD_LOGIC; 
  signal blk00000001_sig0000010a : STD_LOGIC; 
  signal blk00000001_sig00000109 : STD_LOGIC; 
  signal blk00000001_sig00000108 : STD_LOGIC; 
  signal blk00000001_sig00000107 : STD_LOGIC; 
  signal blk00000001_sig00000106 : STD_LOGIC; 
  signal blk00000001_sig00000105 : STD_LOGIC; 
  signal blk00000001_sig00000104 : STD_LOGIC; 
  signal blk00000001_sig00000103 : STD_LOGIC; 
  signal blk00000001_sig00000102 : STD_LOGIC; 
  signal blk00000001_sig00000101 : STD_LOGIC; 
  signal blk00000001_sig00000100 : STD_LOGIC; 
  signal blk00000001_sig000000ff : STD_LOGIC; 
  signal blk00000001_sig000000fe : STD_LOGIC; 
  signal blk00000001_sig000000fd : STD_LOGIC; 
  signal blk00000001_sig000000fc : STD_LOGIC; 
  signal blk00000001_sig000000fb : STD_LOGIC; 
  signal blk00000001_sig000000fa : STD_LOGIC; 
  signal blk00000001_sig000000f9 : STD_LOGIC; 
  signal blk00000001_sig000000f8 : STD_LOGIC; 
  signal blk00000001_sig000000f7 : STD_LOGIC; 
  signal blk00000001_sig000000f6 : STD_LOGIC; 
  signal blk00000001_sig000000f5 : STD_LOGIC; 
  signal blk00000001_sig000000f4 : STD_LOGIC; 
  signal blk00000001_sig000000f3 : STD_LOGIC; 
  signal blk00000001_sig000000f2 : STD_LOGIC; 
  signal blk00000001_sig000000f1 : STD_LOGIC; 
  signal blk00000001_sig000000f0 : STD_LOGIC; 
  signal blk00000001_sig000000ef : STD_LOGIC; 
  signal blk00000001_sig000000ee : STD_LOGIC; 
  signal blk00000001_sig000000ed : STD_LOGIC; 
  signal blk00000001_sig000000ec : STD_LOGIC; 
  signal blk00000001_sig000000eb : STD_LOGIC; 
  signal blk00000001_sig000000ea : STD_LOGIC; 
  signal blk00000001_sig000000e9 : STD_LOGIC; 
  signal blk00000001_sig000000e8 : STD_LOGIC; 
  signal blk00000001_sig000000e7 : STD_LOGIC; 
  signal blk00000001_sig000000e6 : STD_LOGIC; 
  signal blk00000001_sig000000e5 : STD_LOGIC; 
  signal blk00000001_sig000000e4 : STD_LOGIC; 
  signal blk00000001_sig000000e3 : STD_LOGIC; 
  signal blk00000001_sig000000e2 : STD_LOGIC; 
  signal blk00000001_sig000000e1 : STD_LOGIC; 
  signal blk00000001_sig000000e0 : STD_LOGIC; 
  signal blk00000001_sig000000df : STD_LOGIC; 
  signal blk00000001_sig000000de : STD_LOGIC; 
  signal blk00000001_sig000000dd : STD_LOGIC; 
  signal blk00000001_sig000000dc : STD_LOGIC; 
  signal blk00000001_sig000000db : STD_LOGIC; 
  signal blk00000001_sig000000da : STD_LOGIC; 
  signal blk00000001_sig000000d9 : STD_LOGIC; 
  signal blk00000001_sig000000d8 : STD_LOGIC; 
  signal blk00000001_sig000000d7 : STD_LOGIC; 
  signal blk00000001_sig000000d6 : STD_LOGIC; 
  signal blk00000001_sig000000d5 : STD_LOGIC; 
  signal blk00000001_sig000000d4 : STD_LOGIC; 
  signal blk00000001_sig000000d3 : STD_LOGIC; 
  signal blk00000001_sig000000d2 : STD_LOGIC; 
  signal blk00000001_sig000000d1 : STD_LOGIC; 
  signal blk00000001_sig000000d0 : STD_LOGIC; 
  signal blk00000001_sig000000cf : STD_LOGIC; 
  signal blk00000001_sig000000ce : STD_LOGIC; 
  signal blk00000001_sig000000cd : STD_LOGIC; 
  signal blk00000001_sig000000cc : STD_LOGIC; 
  signal blk00000001_sig000000cb : STD_LOGIC; 
  signal blk00000001_sig000000ca : STD_LOGIC; 
  signal blk00000001_sig000000c9 : STD_LOGIC; 
  signal blk00000001_sig000000c8 : STD_LOGIC; 
  signal blk00000001_sig000000c7 : STD_LOGIC; 
  signal blk00000001_sig000000c6 : STD_LOGIC; 
  signal blk00000001_sig000000c5 : STD_LOGIC; 
  signal blk00000001_sig000000c4 : STD_LOGIC; 
  signal blk00000001_sig000000c3 : STD_LOGIC; 
  signal blk00000001_sig000000c2 : STD_LOGIC; 
  signal blk00000001_sig000000c1 : STD_LOGIC; 
  signal blk00000001_sig000000c0 : STD_LOGIC; 
  signal blk00000001_sig000000bf : STD_LOGIC; 
  signal blk00000001_sig000000be : STD_LOGIC; 
  signal blk00000001_sig000000bd : STD_LOGIC; 
  signal blk00000001_sig000000bc : STD_LOGIC; 
  signal blk00000001_sig000000bb : STD_LOGIC; 
  signal blk00000001_sig000000ba : STD_LOGIC; 
  signal blk00000001_sig000000b9 : STD_LOGIC; 
  signal blk00000001_sig000000b8 : STD_LOGIC; 
  signal blk00000001_sig000000b7 : STD_LOGIC; 
  signal blk00000001_sig000000b6 : STD_LOGIC; 
  signal blk00000001_sig000000b5 : STD_LOGIC; 
  signal blk00000001_sig000000b4 : STD_LOGIC; 
  signal blk00000001_sig000000b3 : STD_LOGIC; 
  signal blk00000001_sig000000b2 : STD_LOGIC; 
  signal blk00000001_sig000000b1 : STD_LOGIC; 
  signal blk00000001_sig000000b0 : STD_LOGIC; 
  signal blk00000001_sig000000af : STD_LOGIC; 
  signal blk00000001_sig000000ae : STD_LOGIC; 
  signal blk00000001_sig000000ad : STD_LOGIC; 
  signal blk00000001_sig000000ac : STD_LOGIC; 
  signal blk00000001_sig000000ab : STD_LOGIC; 
  signal blk00000001_sig000000aa : STD_LOGIC; 
  signal blk00000001_sig000000a9 : STD_LOGIC; 
  signal blk00000001_sig000000a8 : STD_LOGIC; 
  signal blk00000001_sig000000a7 : STD_LOGIC; 
  signal blk00000001_sig000000a6 : STD_LOGIC; 
  signal blk00000001_sig000000a5 : STD_LOGIC; 
  signal blk00000001_sig000000a4 : STD_LOGIC; 
  signal blk00000001_sig000000a3 : STD_LOGIC; 
  signal blk00000001_sig000000a2 : STD_LOGIC; 
  signal blk00000001_sig000000a1 : STD_LOGIC; 
  signal blk00000001_sig000000a0 : STD_LOGIC; 
  signal blk00000001_sig0000009f : STD_LOGIC; 
  signal blk00000001_sig0000009e : STD_LOGIC; 
  signal blk00000001_sig0000009d : STD_LOGIC; 
  signal blk00000001_sig0000009c : STD_LOGIC; 
  signal blk00000001_sig0000009b : STD_LOGIC; 
  signal blk00000001_sig0000009a : STD_LOGIC; 
  signal blk00000001_sig00000099 : STD_LOGIC; 
  signal blk00000001_sig00000098 : STD_LOGIC; 
  signal blk00000001_sig00000097 : STD_LOGIC; 
  signal blk00000001_sig00000096 : STD_LOGIC; 
  signal blk00000001_sig00000095 : STD_LOGIC; 
  signal blk00000001_sig00000094 : STD_LOGIC; 
  signal blk00000001_sig00000093 : STD_LOGIC; 
  signal blk00000001_sig00000092 : STD_LOGIC; 
  signal blk00000001_sig00000091 : STD_LOGIC; 
  signal blk00000001_sig00000090 : STD_LOGIC; 
  signal blk00000001_sig0000008f : STD_LOGIC; 
  signal blk00000001_sig0000008e : STD_LOGIC; 
  signal blk00000001_sig0000008d : STD_LOGIC; 
  signal blk00000001_sig0000008c : STD_LOGIC; 
  signal blk00000001_sig0000008b : STD_LOGIC; 
  signal blk00000001_sig0000008a : STD_LOGIC; 
  signal blk00000001_sig0000007d : STD_LOGIC; 
  signal blk00000001_sig0000007c : STD_LOGIC; 
  signal blk00000001_sig0000007b : STD_LOGIC; 
  signal blk00000001_sig0000007a : STD_LOGIC; 
  signal blk00000001_sig00000079 : STD_LOGIC; 
  signal blk00000001_sig00000078 : STD_LOGIC; 
  signal blk00000001_sig00000077 : STD_LOGIC; 
  signal blk00000001_sig00000076 : STD_LOGIC; 
  signal blk00000001_sig00000075 : STD_LOGIC; 
  signal blk00000001_sig00000074 : STD_LOGIC; 
  signal blk00000001_sig00000073 : STD_LOGIC; 
  signal blk00000001_sig00000072 : STD_LOGIC; 
  signal blk00000001_sig00000071 : STD_LOGIC; 
  signal blk00000001_sig00000070 : STD_LOGIC; 
  signal blk00000001_sig0000006f : STD_LOGIC; 
  signal blk00000001_sig0000006e : STD_LOGIC; 
  signal blk00000001_sig0000006d : STD_LOGIC; 
  signal blk00000001_sig0000006c : STD_LOGIC; 
  signal blk00000001_sig0000006b : STD_LOGIC; 
  signal blk00000001_sig0000006a : STD_LOGIC; 
  signal blk00000001_sig00000069 : STD_LOGIC; 
  signal blk00000001_sig00000068 : STD_LOGIC; 
  signal blk00000001_sig00000067 : STD_LOGIC; 
  signal blk00000001_sig00000066 : STD_LOGIC; 
  signal blk00000001_sig00000065 : STD_LOGIC; 
  signal blk00000001_sig00000064 : STD_LOGIC; 
  signal blk00000001_sig00000063 : STD_LOGIC; 
  signal blk00000001_sig00000062 : STD_LOGIC; 
  signal blk00000001_sig00000061 : STD_LOGIC; 
  signal blk00000001_sig00000060 : STD_LOGIC; 
  signal blk00000001_sig0000005f : STD_LOGIC; 
  signal blk00000001_sig0000005e : STD_LOGIC; 
  signal blk00000001_sig0000005d : STD_LOGIC; 
  signal blk00000001_sig0000005c : STD_LOGIC; 
  signal blk00000001_sig0000005b : STD_LOGIC; 
  signal blk00000001_sig0000005a : STD_LOGIC; 
  signal blk00000001_sig00000059 : STD_LOGIC; 
  signal blk00000001_sig00000058 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001005 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001004 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001003 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001002 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001001 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00001000 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fff : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ffe : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ffd : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ffc : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ffb : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ffa : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff9 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff8 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff7 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff6 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff5 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff4 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff3 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff2 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff1 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000ff0 : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fef : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fee : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fed : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fec : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000feb : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fea : STD_LOGIC; 
  signal blk00000001_blk00000025_sig00000fe9 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001086 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001085 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001084 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001083 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001082 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001081 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001080 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107f : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107e : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107d : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107c : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107b : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000107a : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001079 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001078 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001077 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001076 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001075 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001074 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001073 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001072 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001071 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001070 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106f : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106e : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106d : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106c : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106b : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000106a : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001069 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001068 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001067 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001066 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001065 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001064 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001063 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001062 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001061 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001060 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105f : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105e : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105d : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105c : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105b : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000105a : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001059 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001058 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001057 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001056 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001055 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001054 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001052 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001051 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig00001050 : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000104f : STD_LOGIC; 
  signal blk00000001_blk000000b1_sig0000104e : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a8 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a7 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a6 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a5 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a4 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a3 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a2 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a1 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig000010a0 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109f : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109e : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109d : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109c : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109b : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000109a : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001099 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001098 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001097 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001096 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001095 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001092 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001091 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig00001090 : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000108f : STD_LOGIC; 
  signal blk00000001_blk0000010e_sig0000108e : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001142 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001141 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001140 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113f : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113e : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113d : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113c : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113b : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000113a : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001139 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001138 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001137 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001136 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001135 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001134 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001133 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001132 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001131 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001130 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112f : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112e : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112d : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112c : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112b : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000112a : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001129 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001128 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001127 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001126 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001125 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001124 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001123 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001122 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001121 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001120 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111f : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111e : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111d : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111c : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111b : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000111a : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001119 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001118 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001117 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001116 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001115 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001114 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001113 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001112 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001111 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001110 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110f : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110e : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110d : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110c : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110b : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig0000110a : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001109 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001108 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001107 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001106 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001102 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001101 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig00001100 : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig000010ff : STD_LOGIC; 
  signal blk00000001_blk0000012b_sig000010fe : STD_LOGIC; 
  signal blk00000001_blk000007e0_blk000007e1_sig0000114e : STD_LOGIC; 
  signal blk00000001_blk000007e0_blk000007e1_sig0000114d : STD_LOGIC; 
  signal blk00000001_blk000007e0_blk000007e1_sig0000114c : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig000011bb : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000119a : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001199 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001198 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001197 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001196 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001195 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001194 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001193 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001192 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001191 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001190 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118f : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118e : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118d : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118c : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118b : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000118a : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001189 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001188 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001187 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001186 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001185 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001184 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001183 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001182 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001181 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig00001180 : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000117f : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000117e : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000117d : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000117c : STD_LOGIC; 
  signal blk00000001_blk000008e6_sig0000117b : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001228 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001207 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001206 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001205 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001204 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001203 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001202 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001201 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig00001200 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ff : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011fe : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011fd : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011fc : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011fb : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011fa : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f9 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f8 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f7 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f6 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f5 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f4 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f3 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f2 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f1 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011f0 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ef : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ee : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ed : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ec : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011eb : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011ea : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011e9 : STD_LOGIC; 
  signal blk00000001_blk00000909_sig000011e8 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001295 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001274 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001273 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001272 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001271 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001270 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126f : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126e : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126d : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126c : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126b : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000126a : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001269 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001268 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001267 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001266 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001265 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001264 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001263 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001262 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001261 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001260 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125f : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125e : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125d : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125c : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125b : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig0000125a : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001259 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001258 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001257 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001256 : STD_LOGIC; 
  signal blk00000001_blk0000092c_sig00001255 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig00001302 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012e1 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012e0 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012df : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012de : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012dd : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012dc : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012db : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012da : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d9 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d8 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d7 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d6 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d5 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d4 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d3 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d2 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d1 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012d0 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012cf : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012ce : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012cd : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012cc : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012cb : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012ca : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c9 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c8 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c7 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c6 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c5 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c4 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c3 : STD_LOGIC; 
  signal blk00000001_blk0000094f_sig000012c2 : STD_LOGIC; 
  signal blk00000001_blk00000972_blk00000973_sig0000130e : STD_LOGIC; 
  signal blk00000001_blk00000972_blk00000973_sig0000130d : STD_LOGIC; 
  signal blk00000001_blk00000972_blk00000973_sig0000130c : STD_LOGIC; 
  signal blk00000001_blk00000978_blk00000979_sig0000131a : STD_LOGIC; 
  signal blk00000001_blk00000978_blk00000979_sig00001319 : STD_LOGIC; 
  signal blk00000001_blk00000978_blk00000979_sig00001318 : STD_LOGIC; 
  signal blk00000001_blk0000097e_blk0000097f_sig00001326 : STD_LOGIC; 
  signal blk00000001_blk0000097e_blk0000097f_sig00001325 : STD_LOGIC; 
  signal blk00000001_blk0000097e_blk0000097f_sig00001324 : STD_LOGIC; 
  signal blk00000001_blk00000984_blk00000985_sig00001332 : STD_LOGIC; 
  signal blk00000001_blk00000984_blk00000985_sig00001331 : STD_LOGIC; 
  signal blk00000001_blk00000984_blk00000985_sig00001330 : STD_LOGIC; 
  signal blk00000001_blk0000098a_blk0000098b_sig0000133e : STD_LOGIC; 
  signal blk00000001_blk0000098a_blk0000098b_sig0000133d : STD_LOGIC; 
  signal blk00000001_blk0000098a_blk0000098b_sig0000133c : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001356 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001355 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001354 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001353 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001352 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001351 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig00001350 : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig0000134f : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig0000134e : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig0000134d : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig0000134c : STD_LOGIC; 
  signal blk00000001_blk000009c5_sig0000134b : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001366 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001365 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001364 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001363 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001362 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001361 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig00001360 : STD_LOGIC; 
  signal blk00000001_blk000009e2_sig0000135f : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig0000137a : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001379 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001378 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001377 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001376 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001375 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001374 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001373 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001372 : STD_LOGIC; 
  signal blk00000001_blk000009fb_sig00001371 : STD_LOGIC; 
  signal blk00000001_blk00000a0b_blk00000a0c_sig00001385 : STD_LOGIC; 
  signal blk00000001_blk00000a0b_blk00000a0c_sig00001384 : STD_LOGIC; 
  signal blk00000001_blk00000a0b_blk00000a0c_sig00001383 : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig00001391 : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig00001390 : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig0000138f : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig0000138e : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig0000138d : STD_LOGIC; 
  signal blk00000001_blk00000a15_sig0000138c : STD_LOGIC; 
  signal blk00000001_blk00000a1f_blk00000a20_sig000013a5 : STD_LOGIC; 
  signal blk00000001_blk00000a1f_blk00000a20_sig000013a4 : STD_LOGIC; 
  signal blk00000001_blk00000a1f_blk00000a20_sig000013a3 : STD_LOGIC; 
  signal blk00000001_blk00000a25_blk00000a26_sig000013b0 : STD_LOGIC; 
  signal blk00000001_blk00000a25_blk00000a26_sig000013af : STD_LOGIC; 
  signal blk00000001_blk00000a25_blk00000a26_sig000013ae : STD_LOGIC; 
  signal blk00000001_blk00000a2b_blk00000a2c_sig000013bb : STD_LOGIC; 
  signal blk00000001_blk00000a2b_blk00000a2c_sig000013ba : STD_LOGIC; 
  signal blk00000001_blk00000a2b_blk00000a2c_sig000013b9 : STD_LOGIC; 
  signal blk00000001_blk00000a31_blk00000a32_sig000013c6 : STD_LOGIC; 
  signal blk00000001_blk00000a31_blk00000a32_sig000013c5 : STD_LOGIC; 
  signal blk00000001_blk00000a31_blk00000a32_sig000013c4 : STD_LOGIC; 
  signal blk00000001_blk00000a37_blk00000a38_sig000013da : STD_LOGIC; 
  signal blk00000001_blk00000a37_blk00000a38_sig000013d9 : STD_LOGIC; 
  signal blk00000001_blk00000a37_blk00000a38_sig000013d8 : STD_LOGIC; 
  signal blk00000001_blk00000a3d_blk00000a3e_sig000013ee : STD_LOGIC; 
  signal blk00000001_blk00000a3d_blk00000a3e_sig000013ed : STD_LOGIC; 
  signal blk00000001_blk00000a3d_blk00000a3e_sig000013ec : STD_LOGIC; 
  signal blk00000001_blk00000a61_blk00000a62_sig000013fb : STD_LOGIC; 
  signal blk00000001_blk00000a61_blk00000a62_sig000013fa : STD_LOGIC; 
  signal blk00000001_blk00000a61_blk00000a62_sig000013f9 : STD_LOGIC; 
  signal blk00000001_blk00000a67_blk00000a68_sig00001406 : STD_LOGIC; 
  signal blk00000001_blk00000a67_blk00000a68_sig00001405 : STD_LOGIC; 
  signal blk00000001_blk00000a67_blk00000a68_sig00001404 : STD_LOGIC; 
  signal blk00000001_blk00000a6d_blk00000a6e_sig00001413 : STD_LOGIC; 
  signal blk00000001_blk00000a6d_blk00000a6e_sig00001412 : STD_LOGIC; 
  signal blk00000001_blk00000a6d_blk00000a6e_sig00001411 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig0000142d : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig0000142c : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig0000142b : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig0000142a : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001429 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001428 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001427 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001426 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001425 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001424 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001423 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001422 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001421 : STD_LOGIC; 
  signal blk00000001_blk00000a9e_sig00001420 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001447 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001446 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001445 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001444 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001443 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001442 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001441 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig00001440 : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig0000143f : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig0000143e : STD_LOGIC; 
  signal blk00000001_blk00000b3c_sig0000143d : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig00001462 : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig00001461 : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig00001460 : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig0000145f : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig0000145e : STD_LOGIC; 
  signal blk00000001_blk00000b4e_blk00000b4f_sig0000145d : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig0000147d : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig0000147c : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig0000147b : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig0000147a : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig00001479 : STD_LOGIC; 
  signal blk00000001_blk00000b5a_blk00000b5b_sig00001478 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001498 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001497 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001496 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001495 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001494 : STD_LOGIC; 
  signal blk00000001_blk00000b66_blk00000b67_sig00001493 : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014b3 : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014b2 : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014b1 : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014b0 : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014af : STD_LOGIC; 
  signal blk00000001_blk00000b72_blk00000b73_sig000014ae : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d56_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d55_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d54_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d53_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d52_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d51_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d50_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4f_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4e_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4d_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4c_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4b_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d4a_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d49_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d48_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d47_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d46_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d45_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d44_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d43_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d41_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d3f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d3d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d3b_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d39_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d38_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d37_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000d36_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b1b_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b1a_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b0f_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b0d_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b01_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000aff_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000ad3_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000ad1_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000acd_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000acb_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a5e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000611_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000610_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000060f_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000060e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000060d_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000060c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005df_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005de_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005dd_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005dc_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005db_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005da_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005ad_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005ac_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005ab_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005aa_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005a9_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000005a8_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000057b_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000057a_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000579_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000578_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000577_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000576_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000549_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000548_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000547_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000546_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000545_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000544_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000517_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000516_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000515_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000514_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000513_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000512_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e5_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e4_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004e0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004b3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004b2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004b1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004b0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004af_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000004ae_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000043_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000042_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000038_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000037_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000036_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000035_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000025_blk00000034_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk00000103_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk00000102_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000f0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000ef_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000ee_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000ed_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000ec_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000eb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000ea_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000e0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000df_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000de_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000dd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000dc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000db_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000b1_blk000000da_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000010e_blk00000119_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000015d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000015c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000015b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000015a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000159_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000158_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000157_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000156_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000155_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000154_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000153_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000152_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000151_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000150_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000014a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000149_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000148_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000147_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000146_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000145_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000144_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000143_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000142_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000141_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000140_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000013a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000139_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk00000138_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000012e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000012b_blk0000012d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000007e0_blk000007e1_blk000007e4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000008e6_blk00000908_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000008e6_blk00000908_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000008e6_blk00000908_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000008e6_blk00000908_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000909_blk0000092b_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000909_blk0000092b_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000909_blk0000092b_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000909_blk0000092b_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000092c_blk0000094e_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000092c_blk0000094e_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000092c_blk0000094e_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000092c_blk0000094e_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000094f_blk00000971_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000094f_blk00000971_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000094f_blk00000971_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000094f_blk00000971_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000972_blk00000973_blk00000976_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000978_blk00000979_blk0000097c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000097e_blk0000097f_blk00000982_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000984_blk00000985_blk00000988_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk0000098a_blk0000098b_blk0000098e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a0b_blk00000a0c_blk00000a0f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a1f_blk00000a20_blk00000a23_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a25_blk00000a26_blk00000a29_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a2b_blk00000a2c_blk00000a2f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a31_blk00000a32_blk00000a35_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a37_blk00000a38_blk00000a3b_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a3d_blk00000a3e_blk00000a41_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a61_blk00000a62_blk00000a66_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a67_blk00000a68_blk00000a6b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a6d_blk00000a6e_blk00000a72_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000a9e_blk00000aa1_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b58_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b56_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b54_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b52_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b64_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b62_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b60_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b5e_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b66_blk00000b67_blk00000b70_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6e_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6c_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6a_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b72_blk00000b73_blk00000b7c_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b72_blk00000b73_blk00000b7a_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b72_blk00000b73_blk00000b78_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000b72_blk00000b73_blk00000b76_Q31_UNCONNECTED : STD_LOGIC; 
begin
  m_axis_data_tuser(15) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(14) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(13) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(12) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(11) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(10) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(9) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(8) <= NlwRenamedSig_OI_m_axis_data_tuser_8_Q;
  m_axis_data_tuser(7) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(6) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(7) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(6) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(5) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(4) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(3) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(2) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(1) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  s_axis_config_tready <= NlwRenamedSig_OI_s_axis_config_tready;
  s_axis_data_tready <= NlwRenamedSig_OI_s_axis_data_tready;
  m_axis_data_tvalid <= NlwRenamedSig_OI_m_axis_data_tvalid;
  m_axis_status_tvalid <= NlwRenamedSig_OI_m_axis_status_tvalid;
  event_frame_started <= NlwRenamedSig_OI_event_frame_started;
  event_tlast_missing <= NlwRenamedSig_OI_event_tlast_missing;
  event_fft_overflow <= NlwRenamedSig_OI_event_fft_overflow;
  event_status_channel_halt <= NlwRenamedSig_OI_event_status_channel_halt;
  event_data_in_channel_halt <= NlwRenamedSig_OI_event_data_in_channel_halt;
  event_data_out_channel_halt <= NlwRenamedSig_OI_event_data_out_channel_halt;
  blk00000001_blk00000d56 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CEA2 => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d56_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d56_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d56_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d56_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d56_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d56_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(1) => blk00000001_sig000000c0,
      OPMODE(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => blk00000001_sig00000acb,
      C(46) => blk00000001_sig00000acb,
      C(45) => blk00000001_sig00000acb,
      C(44) => blk00000001_sig00000acb,
      C(43) => blk00000001_sig00000aca,
      C(42) => blk00000001_sig00000ac9,
      C(41) => blk00000001_sig00000ac8,
      C(40) => blk00000001_sig00000ac7,
      C(39) => blk00000001_sig00000ac6,
      C(38) => blk00000001_sig00000ac5,
      C(37) => blk00000001_sig00000ac4,
      C(36) => blk00000001_sig00000ac3,
      C(35) => blk00000001_sig00000ac2,
      C(34) => blk00000001_sig00000ac1,
      C(33) => blk00000001_sig00000ac0,
      C(32) => blk00000001_sig00000abf,
      C(31) => blk00000001_sig00000abe,
      C(30) => blk00000001_sig00000abd,
      C(29) => blk00000001_sig00000abc,
      C(28) => blk00000001_sig00000abb,
      C(27) => blk00000001_sig00000aba,
      C(26) => blk00000001_sig00000ab9,
      C(25) => blk00000001_sig00000ab8,
      C(24) => blk00000001_sig00000ab7,
      C(23) => blk00000001_sig00000ae0,
      C(22) => blk00000001_sig00000ae0,
      C(21) => blk00000001_sig00000ae0,
      C(20) => blk00000001_sig00000ae0,
      C(19) => blk00000001_sig00000adf,
      C(18) => blk00000001_sig00000ade,
      C(17) => blk00000001_sig00000add,
      C(16) => blk00000001_sig00000adc,
      C(15) => blk00000001_sig00000adb,
      C(14) => blk00000001_sig00000ada,
      C(13) => blk00000001_sig00000ad9,
      C(12) => blk00000001_sig00000ad8,
      C(11) => blk00000001_sig00000ad7,
      C(10) => blk00000001_sig00000ad6,
      C(9) => blk00000001_sig00000ad5,
      C(8) => blk00000001_sig00000ad4,
      C(7) => blk00000001_sig00000ad3,
      C(6) => blk00000001_sig00000ad2,
      C(5) => blk00000001_sig00000ad1,
      C(4) => blk00000001_sig00000ad0,
      C(3) => blk00000001_sig00000acf,
      C(2) => blk00000001_sig00000ace,
      C(1) => blk00000001_sig00000acd,
      C(0) => blk00000001_sig00000acc,
      B(17) => blk00000001_sig00000a89,
      B(16) => blk00000001_sig00000a88,
      B(15) => blk00000001_sig00000a87,
      B(14) => blk00000001_sig00000a86,
      B(13) => blk00000001_sig00000a85,
      B(12) => blk00000001_sig00000a84,
      B(11) => blk00000001_sig00000a83,
      B(10) => blk00000001_sig00000a82,
      B(9) => blk00000001_sig00000a81,
      B(8) => blk00000001_sig00000a80,
      B(7) => blk00000001_sig00000a7f,
      B(6) => blk00000001_sig00000a7e,
      B(5) => blk00000001_sig00000a7d,
      B(4) => blk00000001_sig00000a7c,
      B(3) => blk00000001_sig00000a7b,
      B(2) => blk00000001_sig00000a7a,
      B(1) => blk00000001_sig00000a79,
      B(0) => blk00000001_sig00000a78,
      P(47) => NLW_blk00000001_blk00000d56_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d56_P_46_UNCONNECTED,
      P(45) => blk00000001_sig00000657,
      P(44) => blk00000001_sig00000656,
      P(43) => blk00000001_sig00000655,
      P(42) => blk00000001_sig00000654,
      P(41) => blk00000001_sig00000653,
      P(40) => blk00000001_sig00000652,
      P(39) => blk00000001_sig00000651,
      P(38) => blk00000001_sig00000650,
      P(37) => blk00000001_sig0000064f,
      P(36) => blk00000001_sig0000064e,
      P(35) => blk00000001_sig0000064d,
      P(34) => blk00000001_sig0000064c,
      P(33) => blk00000001_sig0000064b,
      P(32) => blk00000001_sig0000064a,
      P(31) => blk00000001_sig00000649,
      P(30) => blk00000001_sig00000648,
      P(29) => blk00000001_sig00000647,
      P(28) => blk00000001_sig00000646,
      P(27) => blk00000001_sig00000645,
      P(26) => blk00000001_sig00000644,
      P(25) => blk00000001_sig00000643,
      P(24) => blk00000001_sig00000642,
      P(23) => NLW_blk00000001_blk00000d56_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d56_P_22_UNCONNECTED,
      P(21) => blk00000001_sig0000066d,
      P(20) => blk00000001_sig0000066c,
      P(19) => blk00000001_sig0000066b,
      P(18) => blk00000001_sig0000066a,
      P(17) => blk00000001_sig00000669,
      P(16) => blk00000001_sig00000668,
      P(15) => blk00000001_sig00000667,
      P(14) => blk00000001_sig00000666,
      P(13) => blk00000001_sig00000665,
      P(12) => blk00000001_sig00000664,
      P(11) => blk00000001_sig00000663,
      P(10) => blk00000001_sig00000662,
      P(9) => blk00000001_sig00000661,
      P(8) => blk00000001_sig00000660,
      P(7) => blk00000001_sig0000065f,
      P(6) => blk00000001_sig0000065e,
      P(5) => blk00000001_sig0000065d,
      P(4) => blk00000001_sig0000065c,
      P(3) => blk00000001_sig0000065b,
      P(2) => blk00000001_sig0000065a,
      P(1) => blk00000001_sig00000659,
      P(0) => blk00000001_sig00000658,
      A(29) => blk00000001_sig00000a77,
      A(28) => blk00000001_sig00000a77,
      A(27) => blk00000001_sig00000a77,
      A(26) => blk00000001_sig00000a77,
      A(25) => blk00000001_sig00000a76,
      A(24) => blk00000001_sig00000a75,
      A(23) => blk00000001_sig00000a74,
      A(22) => blk00000001_sig00000a73,
      A(21) => blk00000001_sig00000a72,
      A(20) => blk00000001_sig00000a71,
      A(19) => blk00000001_sig00000a70,
      A(18) => blk00000001_sig00000a6f,
      A(17) => blk00000001_sig00000a6e,
      A(16) => blk00000001_sig00000a6d,
      A(15) => blk00000001_sig00000a6c,
      A(14) => blk00000001_sig00000a6b,
      A(13) => blk00000001_sig00000a6a,
      A(12) => blk00000001_sig00000a69,
      A(11) => blk00000001_sig00000a68,
      A(10) => blk00000001_sig00000a67,
      A(9) => blk00000001_sig00000a66,
      A(8) => blk00000001_sig00000a65,
      A(7) => blk00000001_sig00000a64,
      A(6) => blk00000001_sig00000a63,
      A(5) => blk00000001_sig00000a8c,
      A(4) => blk00000001_sig00000a8c,
      A(3) => blk00000001_sig00000a8c,
      A(2) => blk00000001_sig00000a8c,
      A(1) => blk00000001_sig00000a8b,
      A(0) => blk00000001_sig00000a8a,
      PCOUT(47) => blk00000001_sig00000c89,
      PCOUT(46) => blk00000001_sig00000c88,
      PCOUT(45) => blk00000001_sig00000c87,
      PCOUT(44) => blk00000001_sig00000c86,
      PCOUT(43) => blk00000001_sig00000c85,
      PCOUT(42) => blk00000001_sig00000c84,
      PCOUT(41) => blk00000001_sig00000c83,
      PCOUT(40) => blk00000001_sig00000c82,
      PCOUT(39) => blk00000001_sig00000c81,
      PCOUT(38) => blk00000001_sig00000c80,
      PCOUT(37) => blk00000001_sig00000c7f,
      PCOUT(36) => blk00000001_sig00000c7e,
      PCOUT(35) => blk00000001_sig00000c7d,
      PCOUT(34) => blk00000001_sig00000c7c,
      PCOUT(33) => blk00000001_sig00000c7b,
      PCOUT(32) => blk00000001_sig00000c7a,
      PCOUT(31) => blk00000001_sig00000c79,
      PCOUT(30) => blk00000001_sig00000c78,
      PCOUT(29) => blk00000001_sig00000c77,
      PCOUT(28) => blk00000001_sig00000c76,
      PCOUT(27) => blk00000001_sig00000c75,
      PCOUT(26) => blk00000001_sig00000c74,
      PCOUT(25) => blk00000001_sig00000c73,
      PCOUT(24) => blk00000001_sig00000c72,
      PCOUT(23) => blk00000001_sig00000c71,
      PCOUT(22) => blk00000001_sig00000c70,
      PCOUT(21) => blk00000001_sig00000c6f,
      PCOUT(20) => blk00000001_sig00000c6e,
      PCOUT(19) => blk00000001_sig00000c6d,
      PCOUT(18) => blk00000001_sig00000c6c,
      PCOUT(17) => blk00000001_sig00000c6b,
      PCOUT(16) => blk00000001_sig00000c6a,
      PCOUT(15) => blk00000001_sig00000c69,
      PCOUT(14) => blk00000001_sig00000c68,
      PCOUT(13) => blk00000001_sig00000c67,
      PCOUT(12) => blk00000001_sig00000c66,
      PCOUT(11) => blk00000001_sig00000c65,
      PCOUT(10) => blk00000001_sig00000c64,
      PCOUT(9) => blk00000001_sig00000c63,
      PCOUT(8) => blk00000001_sig00000c62,
      PCOUT(7) => blk00000001_sig00000c61,
      PCOUT(6) => blk00000001_sig00000c60,
      PCOUT(5) => blk00000001_sig00000c5f,
      PCOUT(4) => blk00000001_sig00000c5e,
      PCOUT(3) => blk00000001_sig00000c5d,
      PCOUT(2) => blk00000001_sig00000c5c,
      PCOUT(1) => blk00000001_sig00000c5b,
      PCOUT(0) => blk00000001_sig00000c5a,
      ACOUT(29) => NLW_blk00000001_blk00000d56_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d56_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d56_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d56_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d56_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d56_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d56_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d56_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d56_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d56_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d56_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d56_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d56_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d56_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d56_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d56_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d56_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d56_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d56_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d56_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d56_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d56_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d56_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d56_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d56_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d56_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d56_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d56_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d56_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d56_ACOUT_0_UNCONNECTED,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d56_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d56_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d56_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d56_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d56_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d56_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d56_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d56_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d56_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d56_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d56_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d56_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d56_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d56_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d56_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d56_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d56_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d56_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d56_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d56_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d56_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d56_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d55 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CEA2 => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d55_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d55_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d55_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d55_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d55_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d55_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(1) => blk00000001_sig000000c0,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000c89,
      PCIN(46) => blk00000001_sig00000c88,
      PCIN(45) => blk00000001_sig00000c87,
      PCIN(44) => blk00000001_sig00000c86,
      PCIN(43) => blk00000001_sig00000c85,
      PCIN(42) => blk00000001_sig00000c84,
      PCIN(41) => blk00000001_sig00000c83,
      PCIN(40) => blk00000001_sig00000c82,
      PCIN(39) => blk00000001_sig00000c81,
      PCIN(38) => blk00000001_sig00000c80,
      PCIN(37) => blk00000001_sig00000c7f,
      PCIN(36) => blk00000001_sig00000c7e,
      PCIN(35) => blk00000001_sig00000c7d,
      PCIN(34) => blk00000001_sig00000c7c,
      PCIN(33) => blk00000001_sig00000c7b,
      PCIN(32) => blk00000001_sig00000c7a,
      PCIN(31) => blk00000001_sig00000c79,
      PCIN(30) => blk00000001_sig00000c78,
      PCIN(29) => blk00000001_sig00000c77,
      PCIN(28) => blk00000001_sig00000c76,
      PCIN(27) => blk00000001_sig00000c75,
      PCIN(26) => blk00000001_sig00000c74,
      PCIN(25) => blk00000001_sig00000c73,
      PCIN(24) => blk00000001_sig00000c72,
      PCIN(23) => blk00000001_sig00000c71,
      PCIN(22) => blk00000001_sig00000c70,
      PCIN(21) => blk00000001_sig00000c6f,
      PCIN(20) => blk00000001_sig00000c6e,
      PCIN(19) => blk00000001_sig00000c6d,
      PCIN(18) => blk00000001_sig00000c6c,
      PCIN(17) => blk00000001_sig00000c6b,
      PCIN(16) => blk00000001_sig00000c6a,
      PCIN(15) => blk00000001_sig00000c69,
      PCIN(14) => blk00000001_sig00000c68,
      PCIN(13) => blk00000001_sig00000c67,
      PCIN(12) => blk00000001_sig00000c66,
      PCIN(11) => blk00000001_sig00000c65,
      PCIN(10) => blk00000001_sig00000c64,
      PCIN(9) => blk00000001_sig00000c63,
      PCIN(8) => blk00000001_sig00000c62,
      PCIN(7) => blk00000001_sig00000c61,
      PCIN(6) => blk00000001_sig00000c60,
      PCIN(5) => blk00000001_sig00000c5f,
      PCIN(4) => blk00000001_sig00000c5e,
      PCIN(3) => blk00000001_sig00000c5d,
      PCIN(2) => blk00000001_sig00000c5c,
      PCIN(1) => blk00000001_sig00000c5b,
      PCIN(0) => blk00000001_sig00000c5a,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig000000c0,
      ALUMODE(0) => blk00000001_sig000000c0,
      C(47) => blk00000001_sig00000acb,
      C(46) => blk00000001_sig00000acb,
      C(45) => blk00000001_sig00000acb,
      C(44) => blk00000001_sig00000acb,
      C(43) => blk00000001_sig00000aca,
      C(42) => blk00000001_sig00000ac9,
      C(41) => blk00000001_sig00000ac8,
      C(40) => blk00000001_sig00000ac7,
      C(39) => blk00000001_sig00000ac6,
      C(38) => blk00000001_sig00000ac5,
      C(37) => blk00000001_sig00000ac4,
      C(36) => blk00000001_sig00000ac3,
      C(35) => blk00000001_sig00000ac2,
      C(34) => blk00000001_sig00000ac1,
      C(33) => blk00000001_sig00000ac0,
      C(32) => blk00000001_sig00000abf,
      C(31) => blk00000001_sig00000abe,
      C(30) => blk00000001_sig00000abd,
      C(29) => blk00000001_sig00000abc,
      C(28) => blk00000001_sig00000abb,
      C(27) => blk00000001_sig00000aba,
      C(26) => blk00000001_sig00000ab9,
      C(25) => blk00000001_sig00000ab8,
      C(24) => blk00000001_sig00000ab7,
      C(23) => blk00000001_sig00000ae0,
      C(22) => blk00000001_sig00000ae0,
      C(21) => blk00000001_sig00000ae0,
      C(20) => blk00000001_sig00000ae0,
      C(19) => blk00000001_sig00000adf,
      C(18) => blk00000001_sig00000ade,
      C(17) => blk00000001_sig00000add,
      C(16) => blk00000001_sig00000adc,
      C(15) => blk00000001_sig00000adb,
      C(14) => blk00000001_sig00000ada,
      C(13) => blk00000001_sig00000ad9,
      C(12) => blk00000001_sig00000ad8,
      C(11) => blk00000001_sig00000ad7,
      C(10) => blk00000001_sig00000ad6,
      C(9) => blk00000001_sig00000ad5,
      C(8) => blk00000001_sig00000ad4,
      C(7) => blk00000001_sig00000ad3,
      C(6) => blk00000001_sig00000ad2,
      C(5) => blk00000001_sig00000ad1,
      C(4) => blk00000001_sig00000ad0,
      C(3) => blk00000001_sig00000acf,
      C(2) => blk00000001_sig00000ace,
      C(1) => blk00000001_sig00000acd,
      C(0) => blk00000001_sig00000acc,
      B(17) => blk00000001_sig00000a89,
      B(16) => blk00000001_sig00000a88,
      B(15) => blk00000001_sig00000a87,
      B(14) => blk00000001_sig00000a86,
      B(13) => blk00000001_sig00000a85,
      B(12) => blk00000001_sig00000a84,
      B(11) => blk00000001_sig00000a83,
      B(10) => blk00000001_sig00000a82,
      B(9) => blk00000001_sig00000a81,
      B(8) => blk00000001_sig00000a80,
      B(7) => blk00000001_sig00000a7f,
      B(6) => blk00000001_sig00000a7e,
      B(5) => blk00000001_sig00000a7d,
      B(4) => blk00000001_sig00000a7c,
      B(3) => blk00000001_sig00000a7b,
      B(2) => blk00000001_sig00000a7a,
      B(1) => blk00000001_sig00000a79,
      B(0) => blk00000001_sig00000a78,
      P(47) => NLW_blk00000001_blk00000d55_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d55_P_46_UNCONNECTED,
      P(45) => blk00000001_sig0000062b,
      P(44) => blk00000001_sig0000062a,
      P(43) => blk00000001_sig00000629,
      P(42) => blk00000001_sig00000628,
      P(41) => blk00000001_sig00000627,
      P(40) => blk00000001_sig00000626,
      P(39) => blk00000001_sig00000625,
      P(38) => blk00000001_sig00000624,
      P(37) => blk00000001_sig00000623,
      P(36) => blk00000001_sig00000622,
      P(35) => blk00000001_sig00000621,
      P(34) => blk00000001_sig00000620,
      P(33) => blk00000001_sig0000061f,
      P(32) => blk00000001_sig0000061e,
      P(31) => blk00000001_sig0000061d,
      P(30) => blk00000001_sig0000061c,
      P(29) => blk00000001_sig0000061b,
      P(28) => blk00000001_sig0000061a,
      P(27) => blk00000001_sig00000619,
      P(26) => blk00000001_sig00000618,
      P(25) => blk00000001_sig00000617,
      P(24) => blk00000001_sig00000616,
      P(23) => NLW_blk00000001_blk00000d55_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d55_P_22_UNCONNECTED,
      P(21) => blk00000001_sig00000641,
      P(20) => blk00000001_sig00000640,
      P(19) => blk00000001_sig0000063f,
      P(18) => blk00000001_sig0000063e,
      P(17) => blk00000001_sig0000063d,
      P(16) => blk00000001_sig0000063c,
      P(15) => blk00000001_sig0000063b,
      P(14) => blk00000001_sig0000063a,
      P(13) => blk00000001_sig00000639,
      P(12) => blk00000001_sig00000638,
      P(11) => blk00000001_sig00000637,
      P(10) => blk00000001_sig00000636,
      P(9) => blk00000001_sig00000635,
      P(8) => blk00000001_sig00000634,
      P(7) => blk00000001_sig00000633,
      P(6) => blk00000001_sig00000632,
      P(5) => blk00000001_sig00000631,
      P(4) => blk00000001_sig00000630,
      P(3) => blk00000001_sig0000062f,
      P(2) => blk00000001_sig0000062e,
      P(1) => blk00000001_sig0000062d,
      P(0) => blk00000001_sig0000062c,
      A(29) => blk00000001_sig00000a77,
      A(28) => blk00000001_sig00000a77,
      A(27) => blk00000001_sig00000a77,
      A(26) => blk00000001_sig00000a77,
      A(25) => blk00000001_sig00000a76,
      A(24) => blk00000001_sig00000a75,
      A(23) => blk00000001_sig00000a74,
      A(22) => blk00000001_sig00000a73,
      A(21) => blk00000001_sig00000a72,
      A(20) => blk00000001_sig00000a71,
      A(19) => blk00000001_sig00000a70,
      A(18) => blk00000001_sig00000a6f,
      A(17) => blk00000001_sig00000a6e,
      A(16) => blk00000001_sig00000a6d,
      A(15) => blk00000001_sig00000a6c,
      A(14) => blk00000001_sig00000a6b,
      A(13) => blk00000001_sig00000a6a,
      A(12) => blk00000001_sig00000a69,
      A(11) => blk00000001_sig00000a68,
      A(10) => blk00000001_sig00000a67,
      A(9) => blk00000001_sig00000a66,
      A(8) => blk00000001_sig00000a65,
      A(7) => blk00000001_sig00000a64,
      A(6) => blk00000001_sig00000a63,
      A(5) => blk00000001_sig00000a8c,
      A(4) => blk00000001_sig00000a8c,
      A(3) => blk00000001_sig00000a8c,
      A(2) => blk00000001_sig00000a8c,
      A(1) => blk00000001_sig00000a8b,
      A(0) => blk00000001_sig00000a8a,
      ACOUT(29) => NLW_blk00000001_blk00000d55_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d55_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d55_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d55_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d55_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d55_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d55_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d55_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d55_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d55_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d55_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d55_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d55_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d55_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d55_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d55_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d55_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d55_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d55_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d55_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d55_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d55_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d55_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d55_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d55_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d55_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d55_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d55_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d55_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d55_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000001_blk00000d55_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d55_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d55_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d55_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d55_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d55_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d55_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d55_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d55_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d55_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d55_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d55_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d55_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d55_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d55_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d55_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d55_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d55_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d55_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d55_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d55_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d55_BCOUT_0_UNCONNECTED,
      PCOUT(47) => NLW_blk00000001_blk00000d55_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d55_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d55_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d55_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d55_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d55_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d55_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d55_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d55_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d55_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d55_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d55_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d55_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d55_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d55_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d55_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d55_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d55_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d55_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d55_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d55_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d55_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d55_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d55_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d55_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d55_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d55_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d55_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d55_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d55_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d55_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d55_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d55_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d55_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d55_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d55_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d55_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d55_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d55_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d55_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d55_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d55_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d55_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d55_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d55_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d55_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d55_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d55_PCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d54 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CEA2 => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d54_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d54_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d54_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d54_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d54_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d54_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(1) => blk00000001_sig000000c0,
      OPMODE(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => blk00000001_sig00000af5,
      C(46) => blk00000001_sig00000af5,
      C(45) => blk00000001_sig00000af5,
      C(44) => blk00000001_sig00000af5,
      C(43) => blk00000001_sig00000af4,
      C(42) => blk00000001_sig00000af3,
      C(41) => blk00000001_sig00000af2,
      C(40) => blk00000001_sig00000af1,
      C(39) => blk00000001_sig00000af0,
      C(38) => blk00000001_sig00000aef,
      C(37) => blk00000001_sig00000aee,
      C(36) => blk00000001_sig00000aed,
      C(35) => blk00000001_sig00000aec,
      C(34) => blk00000001_sig00000aeb,
      C(33) => blk00000001_sig00000aea,
      C(32) => blk00000001_sig00000ae9,
      C(31) => blk00000001_sig00000ae8,
      C(30) => blk00000001_sig00000ae7,
      C(29) => blk00000001_sig00000ae6,
      C(28) => blk00000001_sig00000ae5,
      C(27) => blk00000001_sig00000ae4,
      C(26) => blk00000001_sig00000ae3,
      C(25) => blk00000001_sig00000ae2,
      C(24) => blk00000001_sig00000ae1,
      C(23) => blk00000001_sig00000a62,
      C(22) => blk00000001_sig00000a62,
      C(21) => blk00000001_sig00000a62,
      C(20) => blk00000001_sig00000a62,
      C(19) => blk00000001_sig00000a61,
      C(18) => blk00000001_sig00000a60,
      C(17) => blk00000001_sig00000a5f,
      C(16) => blk00000001_sig00000a5e,
      C(15) => blk00000001_sig00000a5d,
      C(14) => blk00000001_sig00000a5c,
      C(13) => blk00000001_sig00000a5b,
      C(12) => blk00000001_sig00000a5a,
      C(11) => blk00000001_sig00000a59,
      C(10) => blk00000001_sig00000a58,
      C(9) => blk00000001_sig00000a57,
      C(8) => blk00000001_sig00000a56,
      C(7) => blk00000001_sig00000a55,
      C(6) => blk00000001_sig00000a54,
      C(5) => blk00000001_sig00000a53,
      C(4) => blk00000001_sig00000a52,
      C(3) => blk00000001_sig00000a51,
      C(2) => blk00000001_sig00000a50,
      C(1) => blk00000001_sig00000a4f,
      C(0) => blk00000001_sig00000a4e,
      B(17) => blk00000001_sig00000ab3,
      B(16) => blk00000001_sig00000ab2,
      B(15) => blk00000001_sig00000ab1,
      B(14) => blk00000001_sig00000ab0,
      B(13) => blk00000001_sig00000aaf,
      B(12) => blk00000001_sig00000aae,
      B(11) => blk00000001_sig00000aad,
      B(10) => blk00000001_sig00000aac,
      B(9) => blk00000001_sig00000aab,
      B(8) => blk00000001_sig00000aaa,
      B(7) => blk00000001_sig00000aa9,
      B(6) => blk00000001_sig00000aa8,
      B(5) => blk00000001_sig00000aa7,
      B(4) => blk00000001_sig00000aa6,
      B(3) => blk00000001_sig00000aa5,
      B(2) => blk00000001_sig00000aa4,
      B(1) => blk00000001_sig00000aa3,
      B(0) => blk00000001_sig00000aa2,
      P(47) => NLW_blk00000001_blk00000d54_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d54_P_46_UNCONNECTED,
      P(45) => blk00000001_sig000006af,
      P(44) => blk00000001_sig000006ae,
      P(43) => blk00000001_sig000006ad,
      P(42) => blk00000001_sig000006ac,
      P(41) => blk00000001_sig000006ab,
      P(40) => blk00000001_sig000006aa,
      P(39) => blk00000001_sig000006a9,
      P(38) => blk00000001_sig000006a8,
      P(37) => blk00000001_sig000006a7,
      P(36) => blk00000001_sig000006a6,
      P(35) => blk00000001_sig000006a5,
      P(34) => blk00000001_sig000006a4,
      P(33) => blk00000001_sig000006a3,
      P(32) => blk00000001_sig000006a2,
      P(31) => blk00000001_sig000006a1,
      P(30) => blk00000001_sig000006a0,
      P(29) => blk00000001_sig0000069f,
      P(28) => blk00000001_sig0000069e,
      P(27) => blk00000001_sig0000069d,
      P(26) => blk00000001_sig0000069c,
      P(25) => blk00000001_sig0000069b,
      P(24) => blk00000001_sig0000069a,
      P(23) => NLW_blk00000001_blk00000d54_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d54_P_22_UNCONNECTED,
      P(21) => blk00000001_sig000006c5,
      P(20) => blk00000001_sig000006c4,
      P(19) => blk00000001_sig000006c3,
      P(18) => blk00000001_sig000006c2,
      P(17) => blk00000001_sig000006c1,
      P(16) => blk00000001_sig000006c0,
      P(15) => blk00000001_sig000006bf,
      P(14) => blk00000001_sig000006be,
      P(13) => blk00000001_sig000006bd,
      P(12) => blk00000001_sig000006bc,
      P(11) => blk00000001_sig000006bb,
      P(10) => blk00000001_sig000006ba,
      P(9) => blk00000001_sig000006b9,
      P(8) => blk00000001_sig000006b8,
      P(7) => blk00000001_sig000006b7,
      P(6) => blk00000001_sig000006b6,
      P(5) => blk00000001_sig000006b5,
      P(4) => blk00000001_sig000006b4,
      P(3) => blk00000001_sig000006b3,
      P(2) => blk00000001_sig000006b2,
      P(1) => blk00000001_sig000006b1,
      P(0) => blk00000001_sig000006b0,
      A(29) => blk00000001_sig00000aa1,
      A(28) => blk00000001_sig00000aa1,
      A(27) => blk00000001_sig00000aa1,
      A(26) => blk00000001_sig00000aa1,
      A(25) => blk00000001_sig00000aa0,
      A(24) => blk00000001_sig00000a9f,
      A(23) => blk00000001_sig00000a9e,
      A(22) => blk00000001_sig00000a9d,
      A(21) => blk00000001_sig00000a9c,
      A(20) => blk00000001_sig00000a9b,
      A(19) => blk00000001_sig00000a9a,
      A(18) => blk00000001_sig00000a99,
      A(17) => blk00000001_sig00000a98,
      A(16) => blk00000001_sig00000a97,
      A(15) => blk00000001_sig00000a96,
      A(14) => blk00000001_sig00000a95,
      A(13) => blk00000001_sig00000a94,
      A(12) => blk00000001_sig00000a93,
      A(11) => blk00000001_sig00000a92,
      A(10) => blk00000001_sig00000a91,
      A(9) => blk00000001_sig00000a90,
      A(8) => blk00000001_sig00000a8f,
      A(7) => blk00000001_sig00000a8e,
      A(6) => blk00000001_sig00000a8d,
      A(5) => blk00000001_sig00000ab6,
      A(4) => blk00000001_sig00000ab6,
      A(3) => blk00000001_sig00000ab6,
      A(2) => blk00000001_sig00000ab6,
      A(1) => blk00000001_sig00000ab5,
      A(0) => blk00000001_sig00000ab4,
      PCOUT(47) => blk00000001_sig00000c59,
      PCOUT(46) => blk00000001_sig00000c58,
      PCOUT(45) => blk00000001_sig00000c57,
      PCOUT(44) => blk00000001_sig00000c56,
      PCOUT(43) => blk00000001_sig00000c55,
      PCOUT(42) => blk00000001_sig00000c54,
      PCOUT(41) => blk00000001_sig00000c53,
      PCOUT(40) => blk00000001_sig00000c52,
      PCOUT(39) => blk00000001_sig00000c51,
      PCOUT(38) => blk00000001_sig00000c50,
      PCOUT(37) => blk00000001_sig00000c4f,
      PCOUT(36) => blk00000001_sig00000c4e,
      PCOUT(35) => blk00000001_sig00000c4d,
      PCOUT(34) => blk00000001_sig00000c4c,
      PCOUT(33) => blk00000001_sig00000c4b,
      PCOUT(32) => blk00000001_sig00000c4a,
      PCOUT(31) => blk00000001_sig00000c49,
      PCOUT(30) => blk00000001_sig00000c48,
      PCOUT(29) => blk00000001_sig00000c47,
      PCOUT(28) => blk00000001_sig00000c46,
      PCOUT(27) => blk00000001_sig00000c45,
      PCOUT(26) => blk00000001_sig00000c44,
      PCOUT(25) => blk00000001_sig00000c43,
      PCOUT(24) => blk00000001_sig00000c42,
      PCOUT(23) => blk00000001_sig00000c41,
      PCOUT(22) => blk00000001_sig00000c40,
      PCOUT(21) => blk00000001_sig00000c3f,
      PCOUT(20) => blk00000001_sig00000c3e,
      PCOUT(19) => blk00000001_sig00000c3d,
      PCOUT(18) => blk00000001_sig00000c3c,
      PCOUT(17) => blk00000001_sig00000c3b,
      PCOUT(16) => blk00000001_sig00000c3a,
      PCOUT(15) => blk00000001_sig00000c39,
      PCOUT(14) => blk00000001_sig00000c38,
      PCOUT(13) => blk00000001_sig00000c37,
      PCOUT(12) => blk00000001_sig00000c36,
      PCOUT(11) => blk00000001_sig00000c35,
      PCOUT(10) => blk00000001_sig00000c34,
      PCOUT(9) => blk00000001_sig00000c33,
      PCOUT(8) => blk00000001_sig00000c32,
      PCOUT(7) => blk00000001_sig00000c31,
      PCOUT(6) => blk00000001_sig00000c30,
      PCOUT(5) => blk00000001_sig00000c2f,
      PCOUT(4) => blk00000001_sig00000c2e,
      PCOUT(3) => blk00000001_sig00000c2d,
      PCOUT(2) => blk00000001_sig00000c2c,
      PCOUT(1) => blk00000001_sig00000c2b,
      PCOUT(0) => blk00000001_sig00000c2a,
      ACOUT(29) => NLW_blk00000001_blk00000d54_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d54_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d54_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d54_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d54_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d54_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d54_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d54_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d54_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d54_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d54_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d54_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d54_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d54_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d54_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d54_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d54_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d54_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d54_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d54_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d54_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d54_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d54_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d54_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d54_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d54_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d54_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d54_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d54_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d54_ACOUT_0_UNCONNECTED,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d54_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d54_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d54_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d54_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d54_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d54_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d54_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d54_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d54_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d54_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d54_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d54_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d54_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d54_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d54_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d54_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d54_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d54_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d54_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d54_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d54_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d54_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d53 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CEA2 => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d53_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d53_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d53_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d53_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d53_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d53_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(1) => blk00000001_sig000000c0,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000c59,
      PCIN(46) => blk00000001_sig00000c58,
      PCIN(45) => blk00000001_sig00000c57,
      PCIN(44) => blk00000001_sig00000c56,
      PCIN(43) => blk00000001_sig00000c55,
      PCIN(42) => blk00000001_sig00000c54,
      PCIN(41) => blk00000001_sig00000c53,
      PCIN(40) => blk00000001_sig00000c52,
      PCIN(39) => blk00000001_sig00000c51,
      PCIN(38) => blk00000001_sig00000c50,
      PCIN(37) => blk00000001_sig00000c4f,
      PCIN(36) => blk00000001_sig00000c4e,
      PCIN(35) => blk00000001_sig00000c4d,
      PCIN(34) => blk00000001_sig00000c4c,
      PCIN(33) => blk00000001_sig00000c4b,
      PCIN(32) => blk00000001_sig00000c4a,
      PCIN(31) => blk00000001_sig00000c49,
      PCIN(30) => blk00000001_sig00000c48,
      PCIN(29) => blk00000001_sig00000c47,
      PCIN(28) => blk00000001_sig00000c46,
      PCIN(27) => blk00000001_sig00000c45,
      PCIN(26) => blk00000001_sig00000c44,
      PCIN(25) => blk00000001_sig00000c43,
      PCIN(24) => blk00000001_sig00000c42,
      PCIN(23) => blk00000001_sig00000c41,
      PCIN(22) => blk00000001_sig00000c40,
      PCIN(21) => blk00000001_sig00000c3f,
      PCIN(20) => blk00000001_sig00000c3e,
      PCIN(19) => blk00000001_sig00000c3d,
      PCIN(18) => blk00000001_sig00000c3c,
      PCIN(17) => blk00000001_sig00000c3b,
      PCIN(16) => blk00000001_sig00000c3a,
      PCIN(15) => blk00000001_sig00000c39,
      PCIN(14) => blk00000001_sig00000c38,
      PCIN(13) => blk00000001_sig00000c37,
      PCIN(12) => blk00000001_sig00000c36,
      PCIN(11) => blk00000001_sig00000c35,
      PCIN(10) => blk00000001_sig00000c34,
      PCIN(9) => blk00000001_sig00000c33,
      PCIN(8) => blk00000001_sig00000c32,
      PCIN(7) => blk00000001_sig00000c31,
      PCIN(6) => blk00000001_sig00000c30,
      PCIN(5) => blk00000001_sig00000c2f,
      PCIN(4) => blk00000001_sig00000c2e,
      PCIN(3) => blk00000001_sig00000c2d,
      PCIN(2) => blk00000001_sig00000c2c,
      PCIN(1) => blk00000001_sig00000c2b,
      PCIN(0) => blk00000001_sig00000c2a,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig000000c0,
      ALUMODE(0) => blk00000001_sig000000c0,
      C(47) => blk00000001_sig00000af5,
      C(46) => blk00000001_sig00000af5,
      C(45) => blk00000001_sig00000af5,
      C(44) => blk00000001_sig00000af5,
      C(43) => blk00000001_sig00000af4,
      C(42) => blk00000001_sig00000af3,
      C(41) => blk00000001_sig00000af2,
      C(40) => blk00000001_sig00000af1,
      C(39) => blk00000001_sig00000af0,
      C(38) => blk00000001_sig00000aef,
      C(37) => blk00000001_sig00000aee,
      C(36) => blk00000001_sig00000aed,
      C(35) => blk00000001_sig00000aec,
      C(34) => blk00000001_sig00000aeb,
      C(33) => blk00000001_sig00000aea,
      C(32) => blk00000001_sig00000ae9,
      C(31) => blk00000001_sig00000ae8,
      C(30) => blk00000001_sig00000ae7,
      C(29) => blk00000001_sig00000ae6,
      C(28) => blk00000001_sig00000ae5,
      C(27) => blk00000001_sig00000ae4,
      C(26) => blk00000001_sig00000ae3,
      C(25) => blk00000001_sig00000ae2,
      C(24) => blk00000001_sig00000ae1,
      C(23) => blk00000001_sig00000a62,
      C(22) => blk00000001_sig00000a62,
      C(21) => blk00000001_sig00000a62,
      C(20) => blk00000001_sig00000a62,
      C(19) => blk00000001_sig00000a61,
      C(18) => blk00000001_sig00000a60,
      C(17) => blk00000001_sig00000a5f,
      C(16) => blk00000001_sig00000a5e,
      C(15) => blk00000001_sig00000a5d,
      C(14) => blk00000001_sig00000a5c,
      C(13) => blk00000001_sig00000a5b,
      C(12) => blk00000001_sig00000a5a,
      C(11) => blk00000001_sig00000a59,
      C(10) => blk00000001_sig00000a58,
      C(9) => blk00000001_sig00000a57,
      C(8) => blk00000001_sig00000a56,
      C(7) => blk00000001_sig00000a55,
      C(6) => blk00000001_sig00000a54,
      C(5) => blk00000001_sig00000a53,
      C(4) => blk00000001_sig00000a52,
      C(3) => blk00000001_sig00000a51,
      C(2) => blk00000001_sig00000a50,
      C(1) => blk00000001_sig00000a4f,
      C(0) => blk00000001_sig00000a4e,
      B(17) => blk00000001_sig00000ab3,
      B(16) => blk00000001_sig00000ab2,
      B(15) => blk00000001_sig00000ab1,
      B(14) => blk00000001_sig00000ab0,
      B(13) => blk00000001_sig00000aaf,
      B(12) => blk00000001_sig00000aae,
      B(11) => blk00000001_sig00000aad,
      B(10) => blk00000001_sig00000aac,
      B(9) => blk00000001_sig00000aab,
      B(8) => blk00000001_sig00000aaa,
      B(7) => blk00000001_sig00000aa9,
      B(6) => blk00000001_sig00000aa8,
      B(5) => blk00000001_sig00000aa7,
      B(4) => blk00000001_sig00000aa6,
      B(3) => blk00000001_sig00000aa5,
      B(2) => blk00000001_sig00000aa4,
      B(1) => blk00000001_sig00000aa3,
      B(0) => blk00000001_sig00000aa2,
      P(47) => NLW_blk00000001_blk00000d53_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d53_P_46_UNCONNECTED,
      P(45) => blk00000001_sig00000683,
      P(44) => blk00000001_sig00000682,
      P(43) => blk00000001_sig00000681,
      P(42) => blk00000001_sig00000680,
      P(41) => blk00000001_sig0000067f,
      P(40) => blk00000001_sig0000067e,
      P(39) => blk00000001_sig0000067d,
      P(38) => blk00000001_sig0000067c,
      P(37) => blk00000001_sig0000067b,
      P(36) => blk00000001_sig0000067a,
      P(35) => blk00000001_sig00000679,
      P(34) => blk00000001_sig00000678,
      P(33) => blk00000001_sig00000677,
      P(32) => blk00000001_sig00000676,
      P(31) => blk00000001_sig00000675,
      P(30) => blk00000001_sig00000674,
      P(29) => blk00000001_sig00000673,
      P(28) => blk00000001_sig00000672,
      P(27) => blk00000001_sig00000671,
      P(26) => blk00000001_sig00000670,
      P(25) => blk00000001_sig0000066f,
      P(24) => blk00000001_sig0000066e,
      P(23) => NLW_blk00000001_blk00000d53_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d53_P_22_UNCONNECTED,
      P(21) => blk00000001_sig00000699,
      P(20) => blk00000001_sig00000698,
      P(19) => blk00000001_sig00000697,
      P(18) => blk00000001_sig00000696,
      P(17) => blk00000001_sig00000695,
      P(16) => blk00000001_sig00000694,
      P(15) => blk00000001_sig00000693,
      P(14) => blk00000001_sig00000692,
      P(13) => blk00000001_sig00000691,
      P(12) => blk00000001_sig00000690,
      P(11) => blk00000001_sig0000068f,
      P(10) => blk00000001_sig0000068e,
      P(9) => blk00000001_sig0000068d,
      P(8) => blk00000001_sig0000068c,
      P(7) => blk00000001_sig0000068b,
      P(6) => blk00000001_sig0000068a,
      P(5) => blk00000001_sig00000689,
      P(4) => blk00000001_sig00000688,
      P(3) => blk00000001_sig00000687,
      P(2) => blk00000001_sig00000686,
      P(1) => blk00000001_sig00000685,
      P(0) => blk00000001_sig00000684,
      A(29) => blk00000001_sig00000aa1,
      A(28) => blk00000001_sig00000aa1,
      A(27) => blk00000001_sig00000aa1,
      A(26) => blk00000001_sig00000aa1,
      A(25) => blk00000001_sig00000aa0,
      A(24) => blk00000001_sig00000a9f,
      A(23) => blk00000001_sig00000a9e,
      A(22) => blk00000001_sig00000a9d,
      A(21) => blk00000001_sig00000a9c,
      A(20) => blk00000001_sig00000a9b,
      A(19) => blk00000001_sig00000a9a,
      A(18) => blk00000001_sig00000a99,
      A(17) => blk00000001_sig00000a98,
      A(16) => blk00000001_sig00000a97,
      A(15) => blk00000001_sig00000a96,
      A(14) => blk00000001_sig00000a95,
      A(13) => blk00000001_sig00000a94,
      A(12) => blk00000001_sig00000a93,
      A(11) => blk00000001_sig00000a92,
      A(10) => blk00000001_sig00000a91,
      A(9) => blk00000001_sig00000a90,
      A(8) => blk00000001_sig00000a8f,
      A(7) => blk00000001_sig00000a8e,
      A(6) => blk00000001_sig00000a8d,
      A(5) => blk00000001_sig00000ab6,
      A(4) => blk00000001_sig00000ab6,
      A(3) => blk00000001_sig00000ab6,
      A(2) => blk00000001_sig00000ab6,
      A(1) => blk00000001_sig00000ab5,
      A(0) => blk00000001_sig00000ab4,
      ACOUT(29) => NLW_blk00000001_blk00000d53_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d53_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d53_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d53_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d53_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d53_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d53_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d53_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d53_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d53_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d53_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d53_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d53_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d53_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d53_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d53_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d53_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d53_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d53_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d53_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d53_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d53_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d53_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d53_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d53_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d53_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d53_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d53_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d53_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d53_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000001_blk00000d53_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d53_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d53_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d53_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d53_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d53_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d53_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d53_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d53_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d53_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d53_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d53_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d53_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d53_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d53_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d53_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d53_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d53_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d53_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d53_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d53_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d53_BCOUT_0_UNCONNECTED,
      PCOUT(47) => NLW_blk00000001_blk00000d53_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d53_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d53_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d53_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d53_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d53_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d53_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d53_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d53_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d53_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d53_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d53_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d53_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d53_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d53_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d53_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d53_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d53_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d53_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d53_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d53_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d53_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d53_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d53_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d53_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d53_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d53_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d53_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d53_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d53_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d53_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d53_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d53_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d53_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d53_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d53_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d53_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d53_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d53_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d53_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d53_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d53_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d53_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d53_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d53_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d53_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d53_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d53_PCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d52 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CECTRL => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d52_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d52_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d52_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d52_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d52_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d52_OVERFLOW_UNCONNECTED,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig00000ba0,
      OPMODE(4) => blk00000001_sig00000ba0,
      OPMODE(3) => blk00000001_sig00000c01,
      OPMODE(2) => blk00000001_sig00000c01,
      OPMODE(1) => blk00000001_sig00000ba0,
      OPMODE(0) => blk00000001_sig00000ba0,
      C(47) => blk00000001_sig00000615,
      C(46) => blk00000001_sig00000615,
      C(45) => blk00000001_sig00000615,
      C(44) => blk00000001_sig00000615,
      C(43) => blk00000001_sig00000615,
      C(42) => blk00000001_sig00000614,
      C(41) => blk00000001_sig00000613,
      C(40) => blk00000001_sig00000612,
      C(39) => blk00000001_sig00000611,
      C(38) => blk00000001_sig00000610,
      C(37) => blk00000001_sig0000060f,
      C(36) => blk00000001_sig0000060e,
      C(35) => blk00000001_sig0000060d,
      C(34) => blk00000001_sig0000060c,
      C(33) => blk00000001_sig0000060b,
      C(32) => blk00000001_sig0000060a,
      C(31) => blk00000001_sig00000609,
      C(30) => blk00000001_sig00000608,
      C(29) => blk00000001_sig00000607,
      C(28) => blk00000001_sig00000606,
      C(27) => blk00000001_sig00000605,
      C(26) => blk00000001_sig00000604,
      C(25) => blk00000001_sig00000603,
      C(24) => blk00000001_sig00000602,
      C(23) => blk00000001_sig00000501,
      C(22) => blk00000001_sig00000501,
      C(21) => blk00000001_sig00000501,
      C(20) => blk00000001_sig00000501,
      C(19) => blk00000001_sig00000501,
      C(18) => blk00000001_sig00000500,
      C(17) => blk00000001_sig000004ff,
      C(16) => blk00000001_sig000004fe,
      C(15) => blk00000001_sig000004fd,
      C(14) => blk00000001_sig000004fc,
      C(13) => blk00000001_sig000004fb,
      C(12) => blk00000001_sig000004fa,
      C(11) => blk00000001_sig000004f9,
      C(10) => blk00000001_sig000004f8,
      C(9) => blk00000001_sig000004f7,
      C(8) => blk00000001_sig000004f6,
      C(7) => blk00000001_sig000004f5,
      C(6) => blk00000001_sig000004f4,
      C(5) => blk00000001_sig000004f3,
      C(4) => blk00000001_sig000004f2,
      C(3) => blk00000001_sig000004f1,
      C(2) => blk00000001_sig000004f0,
      C(1) => blk00000001_sig000004ef,
      C(0) => blk00000001_sig000004ee,
      B(17) => blk00000001_sig000005d7,
      B(16) => blk00000001_sig000005d6,
      B(15) => blk00000001_sig000005d5,
      B(14) => blk00000001_sig000005d4,
      B(13) => blk00000001_sig000005d3,
      B(12) => blk00000001_sig000005d2,
      B(11) => blk00000001_sig000005d1,
      B(10) => blk00000001_sig000005d0,
      B(9) => blk00000001_sig000005cf,
      B(8) => blk00000001_sig000005ce,
      B(7) => blk00000001_sig000005cd,
      B(6) => blk00000001_sig000005cc,
      B(5) => blk00000001_sig000005cb,
      B(4) => blk00000001_sig000005ca,
      B(3) => blk00000001_sig000005c9,
      B(2) => blk00000001_sig000005c8,
      B(1) => blk00000001_sig000005c7,
      B(0) => blk00000001_sig000005c6,
      P(47) => NLW_blk00000001_blk00000d52_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d52_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d52_P_45_UNCONNECTED,
      P(44) => blk00000001_sig00000b34,
      P(43) => blk00000001_sig00000b33,
      P(42) => blk00000001_sig00000b32,
      P(41) => blk00000001_sig00000b31,
      P(40) => blk00000001_sig00000b30,
      P(39) => blk00000001_sig00000b2f,
      P(38) => blk00000001_sig00000b2e,
      P(37) => blk00000001_sig00000b2d,
      P(36) => blk00000001_sig00000b2c,
      P(35) => blk00000001_sig00000b2b,
      P(34) => blk00000001_sig00000b2a,
      P(33) => blk00000001_sig00000b29,
      P(32) => blk00000001_sig00000b28,
      P(31) => blk00000001_sig00000b27,
      P(30) => blk00000001_sig00000b26,
      P(29) => blk00000001_sig00000b25,
      P(28) => blk00000001_sig00000b24,
      P(27) => blk00000001_sig00000b23,
      P(26) => blk00000001_sig00000b22,
      P(25) => blk00000001_sig00000b21,
      P(24) => blk00000001_sig00000b20,
      P(23) => NLW_blk00000001_blk00000d52_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d52_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d52_P_21_UNCONNECTED,
      P(20) => blk00000001_sig00000b49,
      P(19) => blk00000001_sig00000b48,
      P(18) => blk00000001_sig00000b47,
      P(17) => blk00000001_sig00000b46,
      P(16) => blk00000001_sig00000b45,
      P(15) => blk00000001_sig00000b44,
      P(14) => blk00000001_sig00000b43,
      P(13) => blk00000001_sig00000b42,
      P(12) => blk00000001_sig00000b41,
      P(11) => blk00000001_sig00000b40,
      P(10) => blk00000001_sig00000b3f,
      P(9) => blk00000001_sig00000b3e,
      P(8) => blk00000001_sig00000b3d,
      P(7) => blk00000001_sig00000b3c,
      P(6) => blk00000001_sig00000b3b,
      P(5) => blk00000001_sig00000b3a,
      P(4) => blk00000001_sig00000b39,
      P(3) => blk00000001_sig00000b38,
      P(2) => blk00000001_sig00000b37,
      P(1) => blk00000001_sig00000b36,
      P(0) => blk00000001_sig00000b35,
      A(29) => blk00000001_sig000005c5,
      A(28) => blk00000001_sig000005c5,
      A(27) => blk00000001_sig000005c5,
      A(26) => blk00000001_sig000005c5,
      A(25) => blk00000001_sig000005c5,
      A(24) => blk00000001_sig000005c4,
      A(23) => blk00000001_sig000005c3,
      A(22) => blk00000001_sig000005c2,
      A(21) => blk00000001_sig000005c1,
      A(20) => blk00000001_sig000005c0,
      A(19) => blk00000001_sig000005bf,
      A(18) => blk00000001_sig000005be,
      A(17) => blk00000001_sig000005bd,
      A(16) => blk00000001_sig000005bc,
      A(15) => blk00000001_sig000005bb,
      A(14) => blk00000001_sig000005ba,
      A(13) => blk00000001_sig000005b9,
      A(12) => blk00000001_sig000005b8,
      A(11) => blk00000001_sig000005b7,
      A(10) => blk00000001_sig000005b6,
      A(9) => blk00000001_sig000005b5,
      A(8) => blk00000001_sig000005b4,
      A(7) => blk00000001_sig000005b3,
      A(6) => blk00000001_sig000005b2,
      A(5) => blk00000001_sig000005d9,
      A(4) => blk00000001_sig000005d9,
      A(3) => blk00000001_sig000005d9,
      A(2) => blk00000001_sig000005d9,
      A(1) => blk00000001_sig000005d9,
      A(0) => blk00000001_sig000005d8,
      PCOUT(47) => blk00000001_sig00000c00,
      PCOUT(46) => blk00000001_sig00000bff,
      PCOUT(45) => blk00000001_sig00000bfe,
      PCOUT(44) => blk00000001_sig00000bfd,
      PCOUT(43) => blk00000001_sig00000bfc,
      PCOUT(42) => blk00000001_sig00000bfb,
      PCOUT(41) => blk00000001_sig00000bfa,
      PCOUT(40) => blk00000001_sig00000bf9,
      PCOUT(39) => blk00000001_sig00000bf8,
      PCOUT(38) => blk00000001_sig00000bf7,
      PCOUT(37) => blk00000001_sig00000bf6,
      PCOUT(36) => blk00000001_sig00000bf5,
      PCOUT(35) => blk00000001_sig00000bf4,
      PCOUT(34) => blk00000001_sig00000bf3,
      PCOUT(33) => blk00000001_sig00000bf2,
      PCOUT(32) => blk00000001_sig00000bf1,
      PCOUT(31) => blk00000001_sig00000bf0,
      PCOUT(30) => blk00000001_sig00000bef,
      PCOUT(29) => blk00000001_sig00000bee,
      PCOUT(28) => blk00000001_sig00000bed,
      PCOUT(27) => blk00000001_sig00000bec,
      PCOUT(26) => blk00000001_sig00000beb,
      PCOUT(25) => blk00000001_sig00000bea,
      PCOUT(24) => blk00000001_sig00000be9,
      PCOUT(23) => blk00000001_sig00000be8,
      PCOUT(22) => blk00000001_sig00000be7,
      PCOUT(21) => blk00000001_sig00000be6,
      PCOUT(20) => blk00000001_sig00000be5,
      PCOUT(19) => blk00000001_sig00000be4,
      PCOUT(18) => blk00000001_sig00000be3,
      PCOUT(17) => blk00000001_sig00000be2,
      PCOUT(16) => blk00000001_sig00000be1,
      PCOUT(15) => blk00000001_sig00000be0,
      PCOUT(14) => blk00000001_sig00000bdf,
      PCOUT(13) => blk00000001_sig00000bde,
      PCOUT(12) => blk00000001_sig00000bdd,
      PCOUT(11) => blk00000001_sig00000bdc,
      PCOUT(10) => blk00000001_sig00000bdb,
      PCOUT(9) => blk00000001_sig00000bda,
      PCOUT(8) => blk00000001_sig00000bd9,
      PCOUT(7) => blk00000001_sig00000bd8,
      PCOUT(6) => blk00000001_sig00000bd7,
      PCOUT(5) => blk00000001_sig00000bd6,
      PCOUT(4) => blk00000001_sig00000bd5,
      PCOUT(3) => blk00000001_sig00000bd4,
      PCOUT(2) => blk00000001_sig00000bd3,
      PCOUT(1) => blk00000001_sig00000bd2,
      PCOUT(0) => blk00000001_sig00000bd1,
      ACOUT(29) => NLW_blk00000001_blk00000d52_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d52_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d52_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d52_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d52_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d52_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d52_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d52_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d52_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d52_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d52_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d52_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d52_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d52_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d52_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d52_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d52_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d52_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d52_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d52_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d52_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d52_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d52_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d52_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d52_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d52_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d52_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d52_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d52_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d52_ACOUT_0_UNCONNECTED,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d52_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d52_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d52_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d52_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d52_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d52_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d52_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d52_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d52_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d52_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d52_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d52_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d52_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d52_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d52_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d52_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d52_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d52_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d52_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d52_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d52_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d52_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d51 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CECTRL => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d51_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d51_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d51_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d51_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d51_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d51_OVERFLOW_UNCONNECTED,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000ba0,
      ALUMODE(0) => blk00000001_sig00000ba0,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig00000ba0,
      OPMODE(4) => blk00000001_sig00000ba0,
      OPMODE(3) => blk00000001_sig00000c01,
      OPMODE(2) => blk00000001_sig00000c01,
      OPMODE(1) => blk00000001_sig00000ba0,
      OPMODE(0) => blk00000001_sig00000ba0,
      PCIN(47) => blk00000001_sig00000c00,
      PCIN(46) => blk00000001_sig00000bff,
      PCIN(45) => blk00000001_sig00000bfe,
      PCIN(44) => blk00000001_sig00000bfd,
      PCIN(43) => blk00000001_sig00000bfc,
      PCIN(42) => blk00000001_sig00000bfb,
      PCIN(41) => blk00000001_sig00000bfa,
      PCIN(40) => blk00000001_sig00000bf9,
      PCIN(39) => blk00000001_sig00000bf8,
      PCIN(38) => blk00000001_sig00000bf7,
      PCIN(37) => blk00000001_sig00000bf6,
      PCIN(36) => blk00000001_sig00000bf5,
      PCIN(35) => blk00000001_sig00000bf4,
      PCIN(34) => blk00000001_sig00000bf3,
      PCIN(33) => blk00000001_sig00000bf2,
      PCIN(32) => blk00000001_sig00000bf1,
      PCIN(31) => blk00000001_sig00000bf0,
      PCIN(30) => blk00000001_sig00000bef,
      PCIN(29) => blk00000001_sig00000bee,
      PCIN(28) => blk00000001_sig00000bed,
      PCIN(27) => blk00000001_sig00000bec,
      PCIN(26) => blk00000001_sig00000beb,
      PCIN(25) => blk00000001_sig00000bea,
      PCIN(24) => blk00000001_sig00000be9,
      PCIN(23) => blk00000001_sig00000be8,
      PCIN(22) => blk00000001_sig00000be7,
      PCIN(21) => blk00000001_sig00000be6,
      PCIN(20) => blk00000001_sig00000be5,
      PCIN(19) => blk00000001_sig00000be4,
      PCIN(18) => blk00000001_sig00000be3,
      PCIN(17) => blk00000001_sig00000be2,
      PCIN(16) => blk00000001_sig00000be1,
      PCIN(15) => blk00000001_sig00000be0,
      PCIN(14) => blk00000001_sig00000bdf,
      PCIN(13) => blk00000001_sig00000bde,
      PCIN(12) => blk00000001_sig00000bdd,
      PCIN(11) => blk00000001_sig00000bdc,
      PCIN(10) => blk00000001_sig00000bdb,
      PCIN(9) => blk00000001_sig00000bda,
      PCIN(8) => blk00000001_sig00000bd9,
      PCIN(7) => blk00000001_sig00000bd8,
      PCIN(6) => blk00000001_sig00000bd7,
      PCIN(5) => blk00000001_sig00000bd6,
      PCIN(4) => blk00000001_sig00000bd5,
      PCIN(3) => blk00000001_sig00000bd4,
      PCIN(2) => blk00000001_sig00000bd3,
      PCIN(1) => blk00000001_sig00000bd2,
      PCIN(0) => blk00000001_sig00000bd1,
      C(47) => blk00000001_sig00000c15,
      C(46) => blk00000001_sig00000c15,
      C(45) => blk00000001_sig00000c15,
      C(44) => blk00000001_sig00000c15,
      C(43) => blk00000001_sig00000c15,
      C(42) => blk00000001_sig00000c14,
      C(41) => blk00000001_sig00000c13,
      C(40) => blk00000001_sig00000c12,
      C(39) => blk00000001_sig00000c11,
      C(38) => blk00000001_sig00000c10,
      C(37) => blk00000001_sig00000c0f,
      C(36) => blk00000001_sig00000c0e,
      C(35) => blk00000001_sig00000c0d,
      C(34) => blk00000001_sig00000c0c,
      C(33) => blk00000001_sig00000c0b,
      C(32) => blk00000001_sig00000c0a,
      C(31) => blk00000001_sig00000c09,
      C(30) => blk00000001_sig00000c08,
      C(29) => blk00000001_sig00000c07,
      C(28) => blk00000001_sig00000c06,
      C(27) => blk00000001_sig00000c05,
      C(26) => blk00000001_sig00000c04,
      C(25) => blk00000001_sig00000c03,
      C(24) => blk00000001_sig00000c02,
      C(23) => blk00000001_sig00000c29,
      C(22) => blk00000001_sig00000c29,
      C(21) => blk00000001_sig00000c29,
      C(20) => blk00000001_sig00000c29,
      C(19) => blk00000001_sig00000c29,
      C(18) => blk00000001_sig00000c28,
      C(17) => blk00000001_sig00000c27,
      C(16) => blk00000001_sig00000c26,
      C(15) => blk00000001_sig00000c25,
      C(14) => blk00000001_sig00000c24,
      C(13) => blk00000001_sig00000c23,
      C(12) => blk00000001_sig00000c22,
      C(11) => blk00000001_sig00000c21,
      C(10) => blk00000001_sig00000c20,
      C(9) => blk00000001_sig00000c1f,
      C(8) => blk00000001_sig00000c1e,
      C(7) => blk00000001_sig00000c1d,
      C(6) => blk00000001_sig00000c1c,
      C(5) => blk00000001_sig00000c1b,
      C(4) => blk00000001_sig00000c1a,
      C(3) => blk00000001_sig00000c19,
      C(2) => blk00000001_sig00000c18,
      C(1) => blk00000001_sig00000c17,
      C(0) => blk00000001_sig00000c16,
      B(17) => blk00000001_sig000005c3,
      B(16) => blk00000001_sig000005c2,
      B(15) => blk00000001_sig000005c1,
      B(14) => blk00000001_sig000005c0,
      B(13) => blk00000001_sig000005bf,
      B(12) => blk00000001_sig000005be,
      B(11) => blk00000001_sig000005bd,
      B(10) => blk00000001_sig000005bc,
      B(9) => blk00000001_sig000005bb,
      B(8) => blk00000001_sig000005ba,
      B(7) => blk00000001_sig000005b9,
      B(6) => blk00000001_sig000005b8,
      B(5) => blk00000001_sig000005b7,
      B(4) => blk00000001_sig000005b6,
      B(3) => blk00000001_sig000005b5,
      B(2) => blk00000001_sig000005b4,
      B(1) => blk00000001_sig000005b3,
      B(0) => blk00000001_sig000005b2,
      P(47) => NLW_blk00000001_blk00000d51_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d51_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d51_P_45_UNCONNECTED,
      P(44) => blk00000001_sig00000b0a,
      P(43) => blk00000001_sig00000b09,
      P(42) => blk00000001_sig00000b08,
      P(41) => blk00000001_sig00000b07,
      P(40) => blk00000001_sig00000b06,
      P(39) => blk00000001_sig00000b05,
      P(38) => blk00000001_sig00000b04,
      P(37) => blk00000001_sig00000b03,
      P(36) => blk00000001_sig00000b02,
      P(35) => blk00000001_sig00000b01,
      P(34) => blk00000001_sig00000b00,
      P(33) => blk00000001_sig00000aff,
      P(32) => blk00000001_sig00000afe,
      P(31) => blk00000001_sig00000afd,
      P(30) => blk00000001_sig00000afc,
      P(29) => blk00000001_sig00000afb,
      P(28) => blk00000001_sig00000afa,
      P(27) => blk00000001_sig00000af9,
      P(26) => blk00000001_sig00000af8,
      P(25) => blk00000001_sig00000af7,
      P(24) => blk00000001_sig00000af6,
      P(23) => NLW_blk00000001_blk00000d51_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d51_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d51_P_21_UNCONNECTED,
      P(20) => blk00000001_sig00000b1f,
      P(19) => blk00000001_sig00000b1e,
      P(18) => blk00000001_sig00000b1d,
      P(17) => blk00000001_sig00000b1c,
      P(16) => blk00000001_sig00000b1b,
      P(15) => blk00000001_sig00000b1a,
      P(14) => blk00000001_sig00000b19,
      P(13) => blk00000001_sig00000b18,
      P(12) => blk00000001_sig00000b17,
      P(11) => blk00000001_sig00000b16,
      P(10) => blk00000001_sig00000b15,
      P(9) => blk00000001_sig00000b14,
      P(8) => blk00000001_sig00000b13,
      P(7) => blk00000001_sig00000b12,
      P(6) => blk00000001_sig00000b11,
      P(5) => blk00000001_sig00000b10,
      P(4) => blk00000001_sig00000b0f,
      P(3) => blk00000001_sig00000b0e,
      P(2) => blk00000001_sig00000b0d,
      P(1) => blk00000001_sig00000b0c,
      P(0) => blk00000001_sig00000b0b,
      A(29) => blk00000001_sig00000501,
      A(28) => blk00000001_sig00000501,
      A(27) => blk00000001_sig00000501,
      A(26) => blk00000001_sig00000501,
      A(25) => blk00000001_sig00000501,
      A(24) => blk00000001_sig00000500,
      A(23) => blk00000001_sig000004ff,
      A(22) => blk00000001_sig000004fe,
      A(21) => blk00000001_sig000004fd,
      A(20) => blk00000001_sig000004fc,
      A(19) => blk00000001_sig000004fb,
      A(18) => blk00000001_sig000004fa,
      A(17) => blk00000001_sig000004f9,
      A(16) => blk00000001_sig000004f8,
      A(15) => blk00000001_sig000004f7,
      A(14) => blk00000001_sig000004f6,
      A(13) => blk00000001_sig000004f5,
      A(12) => blk00000001_sig000004f4,
      A(11) => blk00000001_sig000004f3,
      A(10) => blk00000001_sig000004f2,
      A(9) => blk00000001_sig000004f1,
      A(8) => blk00000001_sig000004f0,
      A(7) => blk00000001_sig000004ef,
      A(6) => blk00000001_sig000004ee,
      A(5) => blk00000001_sig000005c5,
      A(4) => blk00000001_sig000005c5,
      A(3) => blk00000001_sig000005c5,
      A(2) => blk00000001_sig000005c5,
      A(1) => blk00000001_sig000005c5,
      A(0) => blk00000001_sig000005c4,
      ACOUT(29) => NLW_blk00000001_blk00000d51_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d51_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d51_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d51_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d51_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d51_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d51_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d51_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d51_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d51_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d51_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d51_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d51_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d51_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d51_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d51_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d51_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d51_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d51_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d51_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d51_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d51_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d51_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d51_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d51_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d51_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d51_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d51_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d51_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d51_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000001_blk00000d51_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d51_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d51_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d51_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d51_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d51_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d51_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d51_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d51_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d51_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d51_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d51_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d51_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d51_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d51_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d51_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d51_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d51_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d51_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d51_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d51_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d51_BCOUT_0_UNCONNECTED,
      PCOUT(47) => NLW_blk00000001_blk00000d51_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d51_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d51_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d51_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d51_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d51_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d51_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d51_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d51_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d51_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d51_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d51_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d51_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d51_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d51_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d51_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d51_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d51_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d51_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d51_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d51_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d51_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d51_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d51_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d51_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d51_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d51_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d51_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d51_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d51_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d51_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d51_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d51_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d51_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d51_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d51_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d51_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d51_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d51_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d51_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d51_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d51_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d51_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d51_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d51_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d51_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d51_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d51_PCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d50 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CECTRL => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d50_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d50_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d50_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d50_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d50_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d50_OVERFLOW_UNCONNECTED,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig00000ba0,
      OPMODE(4) => blk00000001_sig00000ba0,
      OPMODE(3) => blk00000001_sig00000b9f,
      OPMODE(2) => blk00000001_sig00000b9f,
      OPMODE(1) => blk00000001_sig00000b9e,
      OPMODE(0) => blk00000001_sig00000b9e,
      C(47) => blk00000001_sig00000765,
      C(46) => blk00000001_sig00000765,
      C(45) => blk00000001_sig00000765,
      C(44) => blk00000001_sig00000765,
      C(43) => blk00000001_sig00000765,
      C(42) => blk00000001_sig00000765,
      C(41) => blk00000001_sig00000764,
      C(40) => blk00000001_sig00000763,
      C(39) => blk00000001_sig00000762,
      C(38) => blk00000001_sig00000761,
      C(37) => blk00000001_sig00000760,
      C(36) => blk00000001_sig0000075f,
      C(35) => blk00000001_sig0000075e,
      C(34) => blk00000001_sig0000075d,
      C(33) => blk00000001_sig0000075c,
      C(32) => blk00000001_sig0000075b,
      C(31) => blk00000001_sig0000075a,
      C(30) => blk00000001_sig00000759,
      C(29) => blk00000001_sig00000758,
      C(28) => blk00000001_sig00000757,
      C(27) => blk00000001_sig00000756,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => blk00000001_sig00000775,
      C(22) => blk00000001_sig00000775,
      C(21) => blk00000001_sig00000775,
      C(20) => blk00000001_sig00000775,
      C(19) => blk00000001_sig00000775,
      C(18) => blk00000001_sig00000775,
      C(17) => blk00000001_sig00000774,
      C(16) => blk00000001_sig00000773,
      C(15) => blk00000001_sig00000772,
      C(14) => blk00000001_sig00000771,
      C(13) => blk00000001_sig00000770,
      C(12) => blk00000001_sig0000076f,
      C(11) => blk00000001_sig0000076e,
      C(10) => blk00000001_sig0000076d,
      C(9) => blk00000001_sig0000076c,
      C(8) => blk00000001_sig0000076b,
      C(7) => blk00000001_sig0000076a,
      C(6) => blk00000001_sig00000769,
      C(5) => blk00000001_sig00000768,
      C(4) => blk00000001_sig00000767,
      C(3) => blk00000001_sig00000766,
      C(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig000005ff,
      B(16) => blk00000001_sig000005fe,
      B(15) => blk00000001_sig000005fd,
      B(14) => blk00000001_sig000005fc,
      B(13) => blk00000001_sig000005fb,
      B(12) => blk00000001_sig000005fa,
      B(11) => blk00000001_sig000005f9,
      B(10) => blk00000001_sig000005f8,
      B(9) => blk00000001_sig000005f7,
      B(8) => blk00000001_sig000005f6,
      B(7) => blk00000001_sig000005f5,
      B(6) => blk00000001_sig000005f4,
      B(5) => blk00000001_sig000005f3,
      B(4) => blk00000001_sig000005f2,
      B(3) => blk00000001_sig000005f1,
      B(2) => blk00000001_sig000005f0,
      B(1) => blk00000001_sig000005ef,
      B(0) => blk00000001_sig000005ee,
      P(47) => NLW_blk00000001_blk00000d50_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d50_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d50_P_45_UNCONNECTED,
      P(44) => blk00000001_sig00000b88,
      P(43) => blk00000001_sig00000b87,
      P(42) => blk00000001_sig00000b86,
      P(41) => blk00000001_sig00000b85,
      P(40) => blk00000001_sig00000b84,
      P(39) => blk00000001_sig00000b83,
      P(38) => blk00000001_sig00000b82,
      P(37) => blk00000001_sig00000b81,
      P(36) => blk00000001_sig00000b80,
      P(35) => blk00000001_sig00000b7f,
      P(34) => blk00000001_sig00000b7e,
      P(33) => blk00000001_sig00000b7d,
      P(32) => blk00000001_sig00000b7c,
      P(31) => blk00000001_sig00000b7b,
      P(30) => blk00000001_sig00000b7a,
      P(29) => blk00000001_sig00000b79,
      P(28) => blk00000001_sig00000b78,
      P(27) => blk00000001_sig00000b77,
      P(26) => blk00000001_sig00000b76,
      P(25) => blk00000001_sig00000b75,
      P(24) => blk00000001_sig00000b74,
      P(23) => NLW_blk00000001_blk00000d50_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d50_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d50_P_21_UNCONNECTED,
      P(20) => blk00000001_sig00000b9d,
      P(19) => blk00000001_sig00000b9c,
      P(18) => blk00000001_sig00000b9b,
      P(17) => blk00000001_sig00000b9a,
      P(16) => blk00000001_sig00000b99,
      P(15) => blk00000001_sig00000b98,
      P(14) => blk00000001_sig00000b97,
      P(13) => blk00000001_sig00000b96,
      P(12) => blk00000001_sig00000b95,
      P(11) => blk00000001_sig00000b94,
      P(10) => blk00000001_sig00000b93,
      P(9) => blk00000001_sig00000b92,
      P(8) => blk00000001_sig00000b91,
      P(7) => blk00000001_sig00000b90,
      P(6) => blk00000001_sig00000b8f,
      P(5) => blk00000001_sig00000b8e,
      P(4) => blk00000001_sig00000b8d,
      P(3) => blk00000001_sig00000b8c,
      P(2) => blk00000001_sig00000b8b,
      P(1) => blk00000001_sig00000b8a,
      P(0) => blk00000001_sig00000b89,
      A(29) => blk00000001_sig000005ed,
      A(28) => blk00000001_sig000005ed,
      A(27) => blk00000001_sig000005ed,
      A(26) => blk00000001_sig000005ed,
      A(25) => blk00000001_sig000005ed,
      A(24) => blk00000001_sig000005ec,
      A(23) => blk00000001_sig000005eb,
      A(22) => blk00000001_sig000005ea,
      A(21) => blk00000001_sig000005e9,
      A(20) => blk00000001_sig000005e8,
      A(19) => blk00000001_sig000005e7,
      A(18) => blk00000001_sig000005e6,
      A(17) => blk00000001_sig000005e5,
      A(16) => blk00000001_sig000005e4,
      A(15) => blk00000001_sig000005e3,
      A(14) => blk00000001_sig000005e2,
      A(13) => blk00000001_sig000005e1,
      A(12) => blk00000001_sig000005e0,
      A(11) => blk00000001_sig000005df,
      A(10) => blk00000001_sig000005de,
      A(9) => blk00000001_sig000005dd,
      A(8) => blk00000001_sig000005dc,
      A(7) => blk00000001_sig000005db,
      A(6) => blk00000001_sig000005da,
      A(5) => blk00000001_sig00000601,
      A(4) => blk00000001_sig00000601,
      A(3) => blk00000001_sig00000601,
      A(2) => blk00000001_sig00000601,
      A(1) => blk00000001_sig00000601,
      A(0) => blk00000001_sig00000600,
      PCOUT(47) => blk00000001_sig00000bd0,
      PCOUT(46) => blk00000001_sig00000bcf,
      PCOUT(45) => blk00000001_sig00000bce,
      PCOUT(44) => blk00000001_sig00000bcd,
      PCOUT(43) => blk00000001_sig00000bcc,
      PCOUT(42) => blk00000001_sig00000bcb,
      PCOUT(41) => blk00000001_sig00000bca,
      PCOUT(40) => blk00000001_sig00000bc9,
      PCOUT(39) => blk00000001_sig00000bc8,
      PCOUT(38) => blk00000001_sig00000bc7,
      PCOUT(37) => blk00000001_sig00000bc6,
      PCOUT(36) => blk00000001_sig00000bc5,
      PCOUT(35) => blk00000001_sig00000bc4,
      PCOUT(34) => blk00000001_sig00000bc3,
      PCOUT(33) => blk00000001_sig00000bc2,
      PCOUT(32) => blk00000001_sig00000bc1,
      PCOUT(31) => blk00000001_sig00000bc0,
      PCOUT(30) => blk00000001_sig00000bbf,
      PCOUT(29) => blk00000001_sig00000bbe,
      PCOUT(28) => blk00000001_sig00000bbd,
      PCOUT(27) => blk00000001_sig00000bbc,
      PCOUT(26) => blk00000001_sig00000bbb,
      PCOUT(25) => blk00000001_sig00000bba,
      PCOUT(24) => blk00000001_sig00000bb9,
      PCOUT(23) => blk00000001_sig00000bb8,
      PCOUT(22) => blk00000001_sig00000bb7,
      PCOUT(21) => blk00000001_sig00000bb6,
      PCOUT(20) => blk00000001_sig00000bb5,
      PCOUT(19) => blk00000001_sig00000bb4,
      PCOUT(18) => blk00000001_sig00000bb3,
      PCOUT(17) => blk00000001_sig00000bb2,
      PCOUT(16) => blk00000001_sig00000bb1,
      PCOUT(15) => blk00000001_sig00000bb0,
      PCOUT(14) => blk00000001_sig00000baf,
      PCOUT(13) => blk00000001_sig00000bae,
      PCOUT(12) => blk00000001_sig00000bad,
      PCOUT(11) => blk00000001_sig00000bac,
      PCOUT(10) => blk00000001_sig00000bab,
      PCOUT(9) => blk00000001_sig00000baa,
      PCOUT(8) => blk00000001_sig00000ba9,
      PCOUT(7) => blk00000001_sig00000ba8,
      PCOUT(6) => blk00000001_sig00000ba7,
      PCOUT(5) => blk00000001_sig00000ba6,
      PCOUT(4) => blk00000001_sig00000ba5,
      PCOUT(3) => blk00000001_sig00000ba4,
      PCOUT(2) => blk00000001_sig00000ba3,
      PCOUT(1) => blk00000001_sig00000ba2,
      PCOUT(0) => blk00000001_sig00000ba1,
      ACOUT(29) => NLW_blk00000001_blk00000d50_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d50_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d50_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d50_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d50_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d50_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d50_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d50_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d50_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d50_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d50_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d50_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d50_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d50_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d50_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d50_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d50_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d50_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d50_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d50_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d50_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d50_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d50_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d50_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d50_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d50_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d50_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d50_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d50_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d50_ACOUT_0_UNCONNECTED,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d50_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d50_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d50_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d50_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d50_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d50_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d50_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d50_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d50_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d50_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d50_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d50_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d50_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d50_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d50_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d50_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d50_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d50_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d50_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d50_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d50_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d50_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4f : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "TWO24"
    )
    port map (
      CECTRL => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4f_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4f_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_sig0000008e,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4f_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4f_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4f_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4f_OVERFLOW_UNCONNECTED,
      CEM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000ba0,
      ALUMODE(0) => blk00000001_sig00000ba0,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig00000ba0,
      OPMODE(4) => blk00000001_sig00000ba0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(1) => blk00000001_sig000000c0,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000bd0,
      PCIN(46) => blk00000001_sig00000bcf,
      PCIN(45) => blk00000001_sig00000bce,
      PCIN(44) => blk00000001_sig00000bcd,
      PCIN(43) => blk00000001_sig00000bcc,
      PCIN(42) => blk00000001_sig00000bcb,
      PCIN(41) => blk00000001_sig00000bca,
      PCIN(40) => blk00000001_sig00000bc9,
      PCIN(39) => blk00000001_sig00000bc8,
      PCIN(38) => blk00000001_sig00000bc7,
      PCIN(37) => blk00000001_sig00000bc6,
      PCIN(36) => blk00000001_sig00000bc5,
      PCIN(35) => blk00000001_sig00000bc4,
      PCIN(34) => blk00000001_sig00000bc3,
      PCIN(33) => blk00000001_sig00000bc2,
      PCIN(32) => blk00000001_sig00000bc1,
      PCIN(31) => blk00000001_sig00000bc0,
      PCIN(30) => blk00000001_sig00000bbf,
      PCIN(29) => blk00000001_sig00000bbe,
      PCIN(28) => blk00000001_sig00000bbd,
      PCIN(27) => blk00000001_sig00000bbc,
      PCIN(26) => blk00000001_sig00000bbb,
      PCIN(25) => blk00000001_sig00000bba,
      PCIN(24) => blk00000001_sig00000bb9,
      PCIN(23) => blk00000001_sig00000bb8,
      PCIN(22) => blk00000001_sig00000bb7,
      PCIN(21) => blk00000001_sig00000bb6,
      PCIN(20) => blk00000001_sig00000bb5,
      PCIN(19) => blk00000001_sig00000bb4,
      PCIN(18) => blk00000001_sig00000bb3,
      PCIN(17) => blk00000001_sig00000bb2,
      PCIN(16) => blk00000001_sig00000bb1,
      PCIN(15) => blk00000001_sig00000bb0,
      PCIN(14) => blk00000001_sig00000baf,
      PCIN(13) => blk00000001_sig00000bae,
      PCIN(12) => blk00000001_sig00000bad,
      PCIN(11) => blk00000001_sig00000bac,
      PCIN(10) => blk00000001_sig00000bab,
      PCIN(9) => blk00000001_sig00000baa,
      PCIN(8) => blk00000001_sig00000ba9,
      PCIN(7) => blk00000001_sig00000ba8,
      PCIN(6) => blk00000001_sig00000ba7,
      PCIN(5) => blk00000001_sig00000ba6,
      PCIN(4) => blk00000001_sig00000ba5,
      PCIN(3) => blk00000001_sig00000ba4,
      PCIN(2) => blk00000001_sig00000ba3,
      PCIN(1) => blk00000001_sig00000ba2,
      PCIN(0) => blk00000001_sig00000ba1,
      C(47) => blk00000001_sig00000765,
      C(46) => blk00000001_sig00000765,
      C(45) => blk00000001_sig00000765,
      C(44) => blk00000001_sig00000765,
      C(43) => blk00000001_sig00000765,
      C(42) => blk00000001_sig00000765,
      C(41) => blk00000001_sig00000764,
      C(40) => blk00000001_sig00000763,
      C(39) => blk00000001_sig00000762,
      C(38) => blk00000001_sig00000761,
      C(37) => blk00000001_sig00000760,
      C(36) => blk00000001_sig0000075f,
      C(35) => blk00000001_sig0000075e,
      C(34) => blk00000001_sig0000075d,
      C(33) => blk00000001_sig0000075c,
      C(32) => blk00000001_sig0000075b,
      C(31) => blk00000001_sig0000075a,
      C(30) => blk00000001_sig00000759,
      C(29) => blk00000001_sig00000758,
      C(28) => blk00000001_sig00000757,
      C(27) => blk00000001_sig00000756,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => blk00000001_sig00000775,
      C(22) => blk00000001_sig00000775,
      C(21) => blk00000001_sig00000775,
      C(20) => blk00000001_sig00000775,
      C(19) => blk00000001_sig00000775,
      C(18) => blk00000001_sig00000775,
      C(17) => blk00000001_sig00000774,
      C(16) => blk00000001_sig00000773,
      C(15) => blk00000001_sig00000772,
      C(14) => blk00000001_sig00000771,
      C(13) => blk00000001_sig00000770,
      C(12) => blk00000001_sig0000076f,
      C(11) => blk00000001_sig0000076e,
      C(10) => blk00000001_sig0000076d,
      C(9) => blk00000001_sig0000076c,
      C(8) => blk00000001_sig0000076b,
      C(7) => blk00000001_sig0000076a,
      C(6) => blk00000001_sig00000769,
      C(5) => blk00000001_sig00000768,
      C(4) => blk00000001_sig00000767,
      C(3) => blk00000001_sig00000766,
      C(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig000005ff,
      B(16) => blk00000001_sig000005fe,
      B(15) => blk00000001_sig000005fd,
      B(14) => blk00000001_sig000005fc,
      B(13) => blk00000001_sig000005fb,
      B(12) => blk00000001_sig000005fa,
      B(11) => blk00000001_sig000005f9,
      B(10) => blk00000001_sig000005f8,
      B(9) => blk00000001_sig000005f7,
      B(8) => blk00000001_sig000005f6,
      B(7) => blk00000001_sig000005f5,
      B(6) => blk00000001_sig000005f4,
      B(5) => blk00000001_sig000005f3,
      B(4) => blk00000001_sig000005f2,
      B(3) => blk00000001_sig000005f1,
      B(2) => blk00000001_sig000005f0,
      B(1) => blk00000001_sig000005ef,
      B(0) => blk00000001_sig000005ee,
      P(47) => NLW_blk00000001_blk00000d4f_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4f_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4f_P_45_UNCONNECTED,
      P(44) => blk00000001_sig00000b5e,
      P(43) => blk00000001_sig00000b5d,
      P(42) => blk00000001_sig00000b5c,
      P(41) => blk00000001_sig00000b5b,
      P(40) => blk00000001_sig00000b5a,
      P(39) => blk00000001_sig00000b59,
      P(38) => blk00000001_sig00000b58,
      P(37) => blk00000001_sig00000b57,
      P(36) => blk00000001_sig00000b56,
      P(35) => blk00000001_sig00000b55,
      P(34) => blk00000001_sig00000b54,
      P(33) => blk00000001_sig00000b53,
      P(32) => blk00000001_sig00000b52,
      P(31) => blk00000001_sig00000b51,
      P(30) => blk00000001_sig00000b50,
      P(29) => blk00000001_sig00000b4f,
      P(28) => blk00000001_sig00000b4e,
      P(27) => blk00000001_sig00000b4d,
      P(26) => blk00000001_sig00000b4c,
      P(25) => blk00000001_sig00000b4b,
      P(24) => blk00000001_sig00000b4a,
      P(23) => NLW_blk00000001_blk00000d4f_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d4f_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d4f_P_21_UNCONNECTED,
      P(20) => blk00000001_sig00000b73,
      P(19) => blk00000001_sig00000b72,
      P(18) => blk00000001_sig00000b71,
      P(17) => blk00000001_sig00000b70,
      P(16) => blk00000001_sig00000b6f,
      P(15) => blk00000001_sig00000b6e,
      P(14) => blk00000001_sig00000b6d,
      P(13) => blk00000001_sig00000b6c,
      P(12) => blk00000001_sig00000b6b,
      P(11) => blk00000001_sig00000b6a,
      P(10) => blk00000001_sig00000b69,
      P(9) => blk00000001_sig00000b68,
      P(8) => blk00000001_sig00000b67,
      P(7) => blk00000001_sig00000b66,
      P(6) => blk00000001_sig00000b65,
      P(5) => blk00000001_sig00000b64,
      P(4) => blk00000001_sig00000b63,
      P(3) => blk00000001_sig00000b62,
      P(2) => blk00000001_sig00000b61,
      P(1) => blk00000001_sig00000b60,
      P(0) => blk00000001_sig00000b5f,
      A(29) => blk00000001_sig000005ed,
      A(28) => blk00000001_sig000005ed,
      A(27) => blk00000001_sig000005ed,
      A(26) => blk00000001_sig000005ed,
      A(25) => blk00000001_sig000005ed,
      A(24) => blk00000001_sig000005ec,
      A(23) => blk00000001_sig000005eb,
      A(22) => blk00000001_sig000005ea,
      A(21) => blk00000001_sig000005e9,
      A(20) => blk00000001_sig000005e8,
      A(19) => blk00000001_sig000005e7,
      A(18) => blk00000001_sig000005e6,
      A(17) => blk00000001_sig000005e5,
      A(16) => blk00000001_sig000005e4,
      A(15) => blk00000001_sig000005e3,
      A(14) => blk00000001_sig000005e2,
      A(13) => blk00000001_sig000005e1,
      A(12) => blk00000001_sig000005e0,
      A(11) => blk00000001_sig000005df,
      A(10) => blk00000001_sig000005de,
      A(9) => blk00000001_sig000005dd,
      A(8) => blk00000001_sig000005dc,
      A(7) => blk00000001_sig000005db,
      A(6) => blk00000001_sig000005da,
      A(5) => blk00000001_sig00000601,
      A(4) => blk00000001_sig00000601,
      A(3) => blk00000001_sig00000601,
      A(2) => blk00000001_sig00000601,
      A(1) => blk00000001_sig00000601,
      A(0) => blk00000001_sig00000600,
      ACOUT(29) => NLW_blk00000001_blk00000d4f_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4f_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4f_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4f_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4f_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4f_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4f_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4f_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4f_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4f_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4f_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4f_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4f_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4f_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4f_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4f_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4f_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4f_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4f_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4f_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4f_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4f_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4f_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4f_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4f_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4f_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4f_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4f_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4f_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4f_ACOUT_0_UNCONNECTED,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4f_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4f_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4f_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4f_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4f_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4f_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4f_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4f_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4f_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4f_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4f_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4f_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4f_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4f_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4f_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4f_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4f_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4f_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4f_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4f_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4f_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4f_BCOUT_0_UNCONNECTED,
      PCOUT(47) => NLW_blk00000001_blk00000d4f_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d4f_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d4f_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d4f_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d4f_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d4f_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d4f_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d4f_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d4f_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d4f_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d4f_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d4f_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d4f_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d4f_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d4f_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d4f_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d4f_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d4f_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d4f_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d4f_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d4f_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d4f_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d4f_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d4f_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d4f_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d4f_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d4f_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d4f_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d4f_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d4f_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d4f_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d4f_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d4f_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d4f_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d4f_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d4f_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d4f_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d4f_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d4f_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d4f_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d4f_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d4f_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d4f_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d4f_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d4f_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d4f_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d4f_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d4f_PCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4e : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4e_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4e_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4e_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4e_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4e_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4e_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000984,
      ALUMODE(0) => blk00000001_sig00000984,
      B(17) => blk00000001_sig000008cf,
      B(16) => blk00000001_sig000008cf,
      B(15) => blk00000001_sig000008cf,
      B(14) => blk00000001_sig000008ce,
      B(13) => blk00000001_sig000008cd,
      B(12) => blk00000001_sig000008cc,
      B(11) => blk00000001_sig000008cb,
      B(10) => blk00000001_sig000008ca,
      B(9) => blk00000001_sig000008c9,
      B(8) => blk00000001_sig000008c8,
      B(7) => blk00000001_sig000008c7,
      B(6) => blk00000001_sig000008c6,
      B(5) => blk00000001_sig000008c5,
      B(4) => blk00000001_sig000008c4,
      B(3) => blk00000001_sig000008c3,
      B(2) => blk00000001_sig000008c2,
      B(1) => blk00000001_sig000008c1,
      B(0) => blk00000001_sig000008c0,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000008e0,
      A(23) => blk00000001_sig000008e0,
      A(22) => blk00000001_sig000008e0,
      A(21) => blk00000001_sig000008e0,
      A(20) => blk00000001_sig000008e0,
      A(19) => blk00000001_sig000008e0,
      A(18) => blk00000001_sig000008e0,
      A(17) => blk00000001_sig000008e0,
      A(16) => blk00000001_sig000008e0,
      A(15) => blk00000001_sig000008df,
      A(14) => blk00000001_sig000008de,
      A(13) => blk00000001_sig000008dd,
      A(12) => blk00000001_sig000008dc,
      A(11) => blk00000001_sig000008db,
      A(10) => blk00000001_sig000008da,
      A(9) => blk00000001_sig000008d9,
      A(8) => blk00000001_sig000008d8,
      A(7) => blk00000001_sig000008d7,
      A(6) => blk00000001_sig000008d6,
      A(5) => blk00000001_sig000008d5,
      A(4) => blk00000001_sig000008d4,
      A(3) => blk00000001_sig000008d3,
      A(2) => blk00000001_sig000008d2,
      A(1) => blk00000001_sig000008d1,
      A(0) => blk00000001_sig000008d0,
      PCOUT(47) => blk00000001_sig00000983,
      PCOUT(46) => blk00000001_sig00000982,
      PCOUT(45) => blk00000001_sig00000981,
      PCOUT(44) => blk00000001_sig00000980,
      PCOUT(43) => blk00000001_sig0000097f,
      PCOUT(42) => blk00000001_sig0000097e,
      PCOUT(41) => blk00000001_sig0000097d,
      PCOUT(40) => blk00000001_sig0000097c,
      PCOUT(39) => blk00000001_sig0000097b,
      PCOUT(38) => blk00000001_sig0000097a,
      PCOUT(37) => blk00000001_sig00000979,
      PCOUT(36) => blk00000001_sig00000978,
      PCOUT(35) => blk00000001_sig00000977,
      PCOUT(34) => blk00000001_sig00000976,
      PCOUT(33) => blk00000001_sig00000975,
      PCOUT(32) => blk00000001_sig00000974,
      PCOUT(31) => blk00000001_sig00000973,
      PCOUT(30) => blk00000001_sig00000972,
      PCOUT(29) => blk00000001_sig00000971,
      PCOUT(28) => blk00000001_sig00000970,
      PCOUT(27) => blk00000001_sig0000096f,
      PCOUT(26) => blk00000001_sig0000096e,
      PCOUT(25) => blk00000001_sig0000096d,
      PCOUT(24) => blk00000001_sig0000096c,
      PCOUT(23) => blk00000001_sig0000096b,
      PCOUT(22) => blk00000001_sig0000096a,
      PCOUT(21) => blk00000001_sig00000969,
      PCOUT(20) => blk00000001_sig00000968,
      PCOUT(19) => blk00000001_sig00000967,
      PCOUT(18) => blk00000001_sig00000966,
      PCOUT(17) => blk00000001_sig00000965,
      PCOUT(16) => blk00000001_sig00000964,
      PCOUT(15) => blk00000001_sig00000963,
      PCOUT(14) => blk00000001_sig00000962,
      PCOUT(13) => blk00000001_sig00000961,
      PCOUT(12) => blk00000001_sig00000960,
      PCOUT(11) => blk00000001_sig0000095f,
      PCOUT(10) => blk00000001_sig0000095e,
      PCOUT(9) => blk00000001_sig0000095d,
      PCOUT(8) => blk00000001_sig0000095c,
      PCOUT(7) => blk00000001_sig0000095b,
      PCOUT(6) => blk00000001_sig0000095a,
      PCOUT(5) => blk00000001_sig00000959,
      PCOUT(4) => blk00000001_sig00000958,
      PCOUT(3) => blk00000001_sig00000957,
      PCOUT(2) => blk00000001_sig00000956,
      PCOUT(1) => blk00000001_sig00000955,
      PCOUT(0) => blk00000001_sig00000954,
      ACOUT(29) => NLW_blk00000001_blk00000d4e_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4e_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4e_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4e_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4e_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4e_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4e_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4e_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4e_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4e_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4e_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4e_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4e_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4e_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4e_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4e_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4e_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4e_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4e_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4e_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4e_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4e_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4e_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4e_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4e_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4e_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4e_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4e_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4e_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4e_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4e_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4e_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4e_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4e_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4e_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4e_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4e_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4e_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4e_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4e_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4e_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4e_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4e_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4e_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4e_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4e_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4e_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4e_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4e_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4e_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4e_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4e_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d4e_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4e_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4e_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d4e_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d4e_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d4e_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d4e_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d4e_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d4e_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d4e_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d4e_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d4e_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d4e_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d4e_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d4e_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d4e_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d4e_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d4e_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d4e_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d4e_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d4e_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d4e_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d4e_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d4e_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d4e_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d4e_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d4e_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d4e_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d4e_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d4e_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d4e_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d4e_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d4e_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d4e_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d4e_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d4e_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d4e_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d4e_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d4e_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d4e_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d4e_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d4e_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d4e_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d4e_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d4e_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d4e_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d4e_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d4e_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4d : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4d_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4d_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4d_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4d_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4d_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4d_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000983,
      PCIN(46) => blk00000001_sig00000982,
      PCIN(45) => blk00000001_sig00000981,
      PCIN(44) => blk00000001_sig00000980,
      PCIN(43) => blk00000001_sig0000097f,
      PCIN(42) => blk00000001_sig0000097e,
      PCIN(41) => blk00000001_sig0000097d,
      PCIN(40) => blk00000001_sig0000097c,
      PCIN(39) => blk00000001_sig0000097b,
      PCIN(38) => blk00000001_sig0000097a,
      PCIN(37) => blk00000001_sig00000979,
      PCIN(36) => blk00000001_sig00000978,
      PCIN(35) => blk00000001_sig00000977,
      PCIN(34) => blk00000001_sig00000976,
      PCIN(33) => blk00000001_sig00000975,
      PCIN(32) => blk00000001_sig00000974,
      PCIN(31) => blk00000001_sig00000973,
      PCIN(30) => blk00000001_sig00000972,
      PCIN(29) => blk00000001_sig00000971,
      PCIN(28) => blk00000001_sig00000970,
      PCIN(27) => blk00000001_sig0000096f,
      PCIN(26) => blk00000001_sig0000096e,
      PCIN(25) => blk00000001_sig0000096d,
      PCIN(24) => blk00000001_sig0000096c,
      PCIN(23) => blk00000001_sig0000096b,
      PCIN(22) => blk00000001_sig0000096a,
      PCIN(21) => blk00000001_sig00000969,
      PCIN(20) => blk00000001_sig00000968,
      PCIN(19) => blk00000001_sig00000967,
      PCIN(18) => blk00000001_sig00000966,
      PCIN(17) => blk00000001_sig00000965,
      PCIN(16) => blk00000001_sig00000964,
      PCIN(15) => blk00000001_sig00000963,
      PCIN(14) => blk00000001_sig00000962,
      PCIN(13) => blk00000001_sig00000961,
      PCIN(12) => blk00000001_sig00000960,
      PCIN(11) => blk00000001_sig0000095f,
      PCIN(10) => blk00000001_sig0000095e,
      PCIN(9) => blk00000001_sig0000095d,
      PCIN(8) => blk00000001_sig0000095c,
      PCIN(7) => blk00000001_sig0000095b,
      PCIN(6) => blk00000001_sig0000095a,
      PCIN(5) => blk00000001_sig00000959,
      PCIN(4) => blk00000001_sig00000958,
      PCIN(3) => blk00000001_sig00000957,
      PCIN(2) => blk00000001_sig00000956,
      PCIN(1) => blk00000001_sig00000955,
      PCIN(0) => blk00000001_sig00000954,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000985,
      ALUMODE(0) => blk00000001_sig00000985,
      B(17) => blk00000001_sig000008bf,
      B(16) => blk00000001_sig000008bf,
      B(15) => blk00000001_sig000008bf,
      B(14) => blk00000001_sig000008be,
      B(13) => blk00000001_sig000008bd,
      B(12) => blk00000001_sig000008bc,
      B(11) => blk00000001_sig000008bb,
      B(10) => blk00000001_sig000008ba,
      B(9) => blk00000001_sig000008b9,
      B(8) => blk00000001_sig000008b8,
      B(7) => blk00000001_sig000008b7,
      B(6) => blk00000001_sig000008b6,
      B(5) => blk00000001_sig000008b5,
      B(4) => blk00000001_sig000008b4,
      B(3) => blk00000001_sig000008b3,
      B(2) => blk00000001_sig000008b2,
      B(1) => blk00000001_sig000008b1,
      B(0) => blk00000001_sig000008b0,
      P(47) => NLW_blk00000001_blk00000d4d_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4d_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4d_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d4d_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d4d_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d4d_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d4d_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d4d_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d4d_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d4d_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d4d_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d4d_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d4d_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d4d_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d4d_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d4d_P_32_UNCONNECTED,
      P(31) => blk00000001_sig000006f1,
      P(30) => blk00000001_sig000006f0,
      P(29) => blk00000001_sig000006ef,
      P(28) => blk00000001_sig000006ee,
      P(27) => blk00000001_sig000006ed,
      P(26) => blk00000001_sig000006ec,
      P(25) => blk00000001_sig000006eb,
      P(24) => blk00000001_sig000006ea,
      P(23) => blk00000001_sig000006e9,
      P(22) => blk00000001_sig000006e8,
      P(21) => blk00000001_sig000006e7,
      P(20) => blk00000001_sig000006e6,
      P(19) => blk00000001_sig000006e5,
      P(18) => blk00000001_sig000006e4,
      P(17) => blk00000001_sig000006e3,
      P(16) => blk00000001_sig000006e2,
      P(15) => blk00000001_sig000006e1,
      P(14) => blk00000001_sig000006e0,
      P(13) => blk00000001_sig000006df,
      P(12) => blk00000001_sig000006de,
      P(11) => NLW_blk00000001_blk00000d4d_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d4d_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d4d_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d4d_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d4d_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d4d_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d4d_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d4d_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d4d_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d4d_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d4d_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d4d_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000008f1,
      A(23) => blk00000001_sig000008f1,
      A(22) => blk00000001_sig000008f1,
      A(21) => blk00000001_sig000008f1,
      A(20) => blk00000001_sig000008f1,
      A(19) => blk00000001_sig000008f1,
      A(18) => blk00000001_sig000008f1,
      A(17) => blk00000001_sig000008f1,
      A(16) => blk00000001_sig000008f1,
      A(15) => blk00000001_sig000008f0,
      A(14) => blk00000001_sig000008ef,
      A(13) => blk00000001_sig000008ee,
      A(12) => blk00000001_sig000008ed,
      A(11) => blk00000001_sig000008ec,
      A(10) => blk00000001_sig000008eb,
      A(9) => blk00000001_sig000008ea,
      A(8) => blk00000001_sig000008e9,
      A(7) => blk00000001_sig000008e8,
      A(6) => blk00000001_sig000008e7,
      A(5) => blk00000001_sig000008e6,
      A(4) => blk00000001_sig000008e5,
      A(3) => blk00000001_sig000008e4,
      A(2) => blk00000001_sig000008e3,
      A(1) => blk00000001_sig000008e2,
      A(0) => blk00000001_sig000008e1,
      PCOUT(47) => NLW_blk00000001_blk00000d4d_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d4d_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d4d_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d4d_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d4d_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d4d_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d4d_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d4d_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d4d_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d4d_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d4d_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d4d_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d4d_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d4d_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d4d_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d4d_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d4d_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d4d_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d4d_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d4d_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d4d_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d4d_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d4d_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d4d_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d4d_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d4d_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d4d_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d4d_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d4d_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d4d_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d4d_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d4d_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d4d_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d4d_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d4d_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d4d_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d4d_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d4d_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d4d_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d4d_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d4d_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d4d_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d4d_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d4d_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d4d_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d4d_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d4d_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d4d_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d4d_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4d_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4d_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4d_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4d_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4d_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4d_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4d_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4d_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4d_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4d_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4d_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4d_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4d_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4d_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4d_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4d_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4d_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4d_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4d_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4d_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4d_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4d_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4d_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4d_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4d_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4d_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4d_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4d_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4d_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4d_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4d_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4d_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4d_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4d_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4d_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4d_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4d_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4d_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4d_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4d_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4d_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4d_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4d_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4d_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4d_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4d_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4d_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4d_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4d_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4d_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4d_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4c : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4c_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4c_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4c_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4c_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4c_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4c_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000922,
      ALUMODE(0) => blk00000001_sig00000922,
      B(17) => blk00000001_sig0000085a,
      B(16) => blk00000001_sig0000085a,
      B(15) => blk00000001_sig0000085a,
      B(14) => blk00000001_sig00000859,
      B(13) => blk00000001_sig00000858,
      B(12) => blk00000001_sig00000857,
      B(11) => blk00000001_sig00000856,
      B(10) => blk00000001_sig00000855,
      B(9) => blk00000001_sig00000854,
      B(8) => blk00000001_sig00000853,
      B(7) => blk00000001_sig00000852,
      B(6) => blk00000001_sig00000851,
      B(5) => blk00000001_sig00000850,
      B(4) => blk00000001_sig0000084f,
      B(3) => blk00000001_sig0000084e,
      B(2) => blk00000001_sig0000084d,
      B(1) => blk00000001_sig0000084c,
      B(0) => blk00000001_sig0000084b,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig0000086b,
      A(23) => blk00000001_sig0000086b,
      A(22) => blk00000001_sig0000086b,
      A(21) => blk00000001_sig0000086b,
      A(20) => blk00000001_sig0000086b,
      A(19) => blk00000001_sig0000086b,
      A(18) => blk00000001_sig0000086b,
      A(17) => blk00000001_sig0000086b,
      A(16) => blk00000001_sig0000086b,
      A(15) => blk00000001_sig0000086a,
      A(14) => blk00000001_sig00000869,
      A(13) => blk00000001_sig00000868,
      A(12) => blk00000001_sig00000867,
      A(11) => blk00000001_sig00000866,
      A(10) => blk00000001_sig00000865,
      A(9) => blk00000001_sig00000864,
      A(8) => blk00000001_sig00000863,
      A(7) => blk00000001_sig00000862,
      A(6) => blk00000001_sig00000861,
      A(5) => blk00000001_sig00000860,
      A(4) => blk00000001_sig0000085f,
      A(3) => blk00000001_sig0000085e,
      A(2) => blk00000001_sig0000085d,
      A(1) => blk00000001_sig0000085c,
      A(0) => blk00000001_sig0000085b,
      PCOUT(47) => blk00000001_sig00000953,
      PCOUT(46) => blk00000001_sig00000952,
      PCOUT(45) => blk00000001_sig00000951,
      PCOUT(44) => blk00000001_sig00000950,
      PCOUT(43) => blk00000001_sig0000094f,
      PCOUT(42) => blk00000001_sig0000094e,
      PCOUT(41) => blk00000001_sig0000094d,
      PCOUT(40) => blk00000001_sig0000094c,
      PCOUT(39) => blk00000001_sig0000094b,
      PCOUT(38) => blk00000001_sig0000094a,
      PCOUT(37) => blk00000001_sig00000949,
      PCOUT(36) => blk00000001_sig00000948,
      PCOUT(35) => blk00000001_sig00000947,
      PCOUT(34) => blk00000001_sig00000946,
      PCOUT(33) => blk00000001_sig00000945,
      PCOUT(32) => blk00000001_sig00000944,
      PCOUT(31) => blk00000001_sig00000943,
      PCOUT(30) => blk00000001_sig00000942,
      PCOUT(29) => blk00000001_sig00000941,
      PCOUT(28) => blk00000001_sig00000940,
      PCOUT(27) => blk00000001_sig0000093f,
      PCOUT(26) => blk00000001_sig0000093e,
      PCOUT(25) => blk00000001_sig0000093d,
      PCOUT(24) => blk00000001_sig0000093c,
      PCOUT(23) => blk00000001_sig0000093b,
      PCOUT(22) => blk00000001_sig0000093a,
      PCOUT(21) => blk00000001_sig00000939,
      PCOUT(20) => blk00000001_sig00000938,
      PCOUT(19) => blk00000001_sig00000937,
      PCOUT(18) => blk00000001_sig00000936,
      PCOUT(17) => blk00000001_sig00000935,
      PCOUT(16) => blk00000001_sig00000934,
      PCOUT(15) => blk00000001_sig00000933,
      PCOUT(14) => blk00000001_sig00000932,
      PCOUT(13) => blk00000001_sig00000931,
      PCOUT(12) => blk00000001_sig00000930,
      PCOUT(11) => blk00000001_sig0000092f,
      PCOUT(10) => blk00000001_sig0000092e,
      PCOUT(9) => blk00000001_sig0000092d,
      PCOUT(8) => blk00000001_sig0000092c,
      PCOUT(7) => blk00000001_sig0000092b,
      PCOUT(6) => blk00000001_sig0000092a,
      PCOUT(5) => blk00000001_sig00000929,
      PCOUT(4) => blk00000001_sig00000928,
      PCOUT(3) => blk00000001_sig00000927,
      PCOUT(2) => blk00000001_sig00000926,
      PCOUT(1) => blk00000001_sig00000925,
      PCOUT(0) => blk00000001_sig00000924,
      ACOUT(29) => NLW_blk00000001_blk00000d4c_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4c_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4c_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4c_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4c_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4c_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4c_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4c_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4c_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4c_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4c_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4c_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4c_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4c_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4c_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4c_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4c_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4c_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4c_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4c_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4c_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4c_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4c_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4c_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4c_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4c_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4c_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4c_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4c_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4c_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4c_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4c_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4c_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4c_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4c_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4c_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4c_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4c_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4c_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4c_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4c_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4c_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4c_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4c_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4c_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4c_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4c_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4c_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4c_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4c_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4c_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4c_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d4c_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4c_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4c_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d4c_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d4c_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d4c_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d4c_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d4c_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d4c_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d4c_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d4c_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d4c_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d4c_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d4c_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d4c_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d4c_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d4c_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d4c_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d4c_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d4c_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d4c_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d4c_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d4c_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d4c_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d4c_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d4c_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d4c_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d4c_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d4c_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d4c_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d4c_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d4c_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d4c_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d4c_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d4c_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d4c_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d4c_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d4c_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d4c_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d4c_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d4c_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d4c_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d4c_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d4c_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d4c_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d4c_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d4c_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d4c_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4b : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4b_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4b_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4b_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4b_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4b_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4b_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000953,
      PCIN(46) => blk00000001_sig00000952,
      PCIN(45) => blk00000001_sig00000951,
      PCIN(44) => blk00000001_sig00000950,
      PCIN(43) => blk00000001_sig0000094f,
      PCIN(42) => blk00000001_sig0000094e,
      PCIN(41) => blk00000001_sig0000094d,
      PCIN(40) => blk00000001_sig0000094c,
      PCIN(39) => blk00000001_sig0000094b,
      PCIN(38) => blk00000001_sig0000094a,
      PCIN(37) => blk00000001_sig00000949,
      PCIN(36) => blk00000001_sig00000948,
      PCIN(35) => blk00000001_sig00000947,
      PCIN(34) => blk00000001_sig00000946,
      PCIN(33) => blk00000001_sig00000945,
      PCIN(32) => blk00000001_sig00000944,
      PCIN(31) => blk00000001_sig00000943,
      PCIN(30) => blk00000001_sig00000942,
      PCIN(29) => blk00000001_sig00000941,
      PCIN(28) => blk00000001_sig00000940,
      PCIN(27) => blk00000001_sig0000093f,
      PCIN(26) => blk00000001_sig0000093e,
      PCIN(25) => blk00000001_sig0000093d,
      PCIN(24) => blk00000001_sig0000093c,
      PCIN(23) => blk00000001_sig0000093b,
      PCIN(22) => blk00000001_sig0000093a,
      PCIN(21) => blk00000001_sig00000939,
      PCIN(20) => blk00000001_sig00000938,
      PCIN(19) => blk00000001_sig00000937,
      PCIN(18) => blk00000001_sig00000936,
      PCIN(17) => blk00000001_sig00000935,
      PCIN(16) => blk00000001_sig00000934,
      PCIN(15) => blk00000001_sig00000933,
      PCIN(14) => blk00000001_sig00000932,
      PCIN(13) => blk00000001_sig00000931,
      PCIN(12) => blk00000001_sig00000930,
      PCIN(11) => blk00000001_sig0000092f,
      PCIN(10) => blk00000001_sig0000092e,
      PCIN(9) => blk00000001_sig0000092d,
      PCIN(8) => blk00000001_sig0000092c,
      PCIN(7) => blk00000001_sig0000092b,
      PCIN(6) => blk00000001_sig0000092a,
      PCIN(5) => blk00000001_sig00000929,
      PCIN(4) => blk00000001_sig00000928,
      PCIN(3) => blk00000001_sig00000927,
      PCIN(2) => blk00000001_sig00000926,
      PCIN(1) => blk00000001_sig00000925,
      PCIN(0) => blk00000001_sig00000924,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig0000084a,
      B(16) => blk00000001_sig0000084a,
      B(15) => blk00000001_sig0000084a,
      B(14) => blk00000001_sig00000849,
      B(13) => blk00000001_sig00000848,
      B(12) => blk00000001_sig00000847,
      B(11) => blk00000001_sig00000846,
      B(10) => blk00000001_sig00000845,
      B(9) => blk00000001_sig00000844,
      B(8) => blk00000001_sig00000843,
      B(7) => blk00000001_sig00000842,
      B(6) => blk00000001_sig00000841,
      B(5) => blk00000001_sig00000840,
      B(4) => blk00000001_sig0000083f,
      B(3) => blk00000001_sig0000083e,
      B(2) => blk00000001_sig0000083d,
      B(1) => blk00000001_sig0000083c,
      B(0) => blk00000001_sig0000083b,
      P(47) => NLW_blk00000001_blk00000d4b_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4b_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4b_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d4b_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d4b_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d4b_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d4b_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d4b_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d4b_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d4b_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d4b_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d4b_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d4b_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d4b_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d4b_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d4b_P_32_UNCONNECTED,
      P(31) => blk00000001_sig00000719,
      P(30) => blk00000001_sig00000718,
      P(29) => blk00000001_sig00000717,
      P(28) => blk00000001_sig00000716,
      P(27) => blk00000001_sig00000715,
      P(26) => blk00000001_sig00000714,
      P(25) => blk00000001_sig00000713,
      P(24) => blk00000001_sig00000712,
      P(23) => blk00000001_sig00000711,
      P(22) => blk00000001_sig00000710,
      P(21) => blk00000001_sig0000070f,
      P(20) => blk00000001_sig0000070e,
      P(19) => blk00000001_sig0000070d,
      P(18) => blk00000001_sig0000070c,
      P(17) => blk00000001_sig0000070b,
      P(16) => blk00000001_sig0000070a,
      P(15) => blk00000001_sig00000709,
      P(14) => blk00000001_sig00000708,
      P(13) => blk00000001_sig00000707,
      P(12) => blk00000001_sig00000706,
      P(11) => NLW_blk00000001_blk00000d4b_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d4b_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d4b_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d4b_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d4b_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d4b_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d4b_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d4b_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d4b_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d4b_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d4b_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d4b_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig0000087c,
      A(23) => blk00000001_sig0000087c,
      A(22) => blk00000001_sig0000087c,
      A(21) => blk00000001_sig0000087c,
      A(20) => blk00000001_sig0000087c,
      A(19) => blk00000001_sig0000087c,
      A(18) => blk00000001_sig0000087c,
      A(17) => blk00000001_sig0000087c,
      A(16) => blk00000001_sig0000087c,
      A(15) => blk00000001_sig0000087b,
      A(14) => blk00000001_sig0000087a,
      A(13) => blk00000001_sig00000879,
      A(12) => blk00000001_sig00000878,
      A(11) => blk00000001_sig00000877,
      A(10) => blk00000001_sig00000876,
      A(9) => blk00000001_sig00000875,
      A(8) => blk00000001_sig00000874,
      A(7) => blk00000001_sig00000873,
      A(6) => blk00000001_sig00000872,
      A(5) => blk00000001_sig00000871,
      A(4) => blk00000001_sig00000870,
      A(3) => blk00000001_sig0000086f,
      A(2) => blk00000001_sig0000086e,
      A(1) => blk00000001_sig0000086d,
      A(0) => blk00000001_sig0000086c,
      PCOUT(47) => NLW_blk00000001_blk00000d4b_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d4b_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d4b_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d4b_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d4b_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d4b_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d4b_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d4b_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d4b_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d4b_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d4b_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d4b_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d4b_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d4b_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d4b_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d4b_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d4b_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d4b_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d4b_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d4b_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d4b_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d4b_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d4b_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d4b_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d4b_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d4b_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d4b_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d4b_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d4b_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d4b_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d4b_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d4b_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d4b_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d4b_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d4b_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d4b_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d4b_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d4b_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d4b_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d4b_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d4b_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d4b_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d4b_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d4b_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d4b_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d4b_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d4b_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d4b_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d4b_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4b_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4b_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4b_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4b_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4b_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4b_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4b_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4b_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4b_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4b_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4b_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4b_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4b_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4b_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4b_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4b_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4b_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4b_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4b_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4b_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4b_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4b_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4b_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4b_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4b_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4b_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4b_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4b_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4b_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4b_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4b_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4b_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4b_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4b_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4b_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4b_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4b_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4b_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4b_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4b_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4b_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4b_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4b_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4b_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4b_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4b_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4b_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4b_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4b_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4b_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4b_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d4a : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d4a_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d4a_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d4a_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d4a_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d4a_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d4a_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000922,
      ALUMODE(0) => blk00000001_sig00000922,
      B(17) => blk00000001_sig000007e7,
      B(16) => blk00000001_sig000007e7,
      B(15) => blk00000001_sig000007e7,
      B(14) => blk00000001_sig000007e6,
      B(13) => blk00000001_sig000007e5,
      B(12) => blk00000001_sig000007e4,
      B(11) => blk00000001_sig000007e3,
      B(10) => blk00000001_sig000007e2,
      B(9) => blk00000001_sig000007e1,
      B(8) => blk00000001_sig000007e0,
      B(7) => blk00000001_sig000007df,
      B(6) => blk00000001_sig000007de,
      B(5) => blk00000001_sig000007dd,
      B(4) => blk00000001_sig000007dc,
      B(3) => blk00000001_sig000007db,
      B(2) => blk00000001_sig000007da,
      B(1) => blk00000001_sig000007d9,
      B(0) => blk00000001_sig000007d8,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000007f8,
      A(23) => blk00000001_sig000007f8,
      A(22) => blk00000001_sig000007f8,
      A(21) => blk00000001_sig000007f8,
      A(20) => blk00000001_sig000007f8,
      A(19) => blk00000001_sig000007f8,
      A(18) => blk00000001_sig000007f8,
      A(17) => blk00000001_sig000007f8,
      A(16) => blk00000001_sig000007f8,
      A(15) => blk00000001_sig000007f7,
      A(14) => blk00000001_sig000007f6,
      A(13) => blk00000001_sig000007f5,
      A(12) => blk00000001_sig000007f4,
      A(11) => blk00000001_sig000007f3,
      A(10) => blk00000001_sig000007f2,
      A(9) => blk00000001_sig000007f1,
      A(8) => blk00000001_sig000007f0,
      A(7) => blk00000001_sig000007ef,
      A(6) => blk00000001_sig000007ee,
      A(5) => blk00000001_sig000007ed,
      A(4) => blk00000001_sig000007ec,
      A(3) => blk00000001_sig000007eb,
      A(2) => blk00000001_sig000007ea,
      A(1) => blk00000001_sig000007e9,
      A(0) => blk00000001_sig000007e8,
      PCOUT(47) => blk00000001_sig00000921,
      PCOUT(46) => blk00000001_sig00000920,
      PCOUT(45) => blk00000001_sig0000091f,
      PCOUT(44) => blk00000001_sig0000091e,
      PCOUT(43) => blk00000001_sig0000091d,
      PCOUT(42) => blk00000001_sig0000091c,
      PCOUT(41) => blk00000001_sig0000091b,
      PCOUT(40) => blk00000001_sig0000091a,
      PCOUT(39) => blk00000001_sig00000919,
      PCOUT(38) => blk00000001_sig00000918,
      PCOUT(37) => blk00000001_sig00000917,
      PCOUT(36) => blk00000001_sig00000916,
      PCOUT(35) => blk00000001_sig00000915,
      PCOUT(34) => blk00000001_sig00000914,
      PCOUT(33) => blk00000001_sig00000913,
      PCOUT(32) => blk00000001_sig00000912,
      PCOUT(31) => blk00000001_sig00000911,
      PCOUT(30) => blk00000001_sig00000910,
      PCOUT(29) => blk00000001_sig0000090f,
      PCOUT(28) => blk00000001_sig0000090e,
      PCOUT(27) => blk00000001_sig0000090d,
      PCOUT(26) => blk00000001_sig0000090c,
      PCOUT(25) => blk00000001_sig0000090b,
      PCOUT(24) => blk00000001_sig0000090a,
      PCOUT(23) => blk00000001_sig00000909,
      PCOUT(22) => blk00000001_sig00000908,
      PCOUT(21) => blk00000001_sig00000907,
      PCOUT(20) => blk00000001_sig00000906,
      PCOUT(19) => blk00000001_sig00000905,
      PCOUT(18) => blk00000001_sig00000904,
      PCOUT(17) => blk00000001_sig00000903,
      PCOUT(16) => blk00000001_sig00000902,
      PCOUT(15) => blk00000001_sig00000901,
      PCOUT(14) => blk00000001_sig00000900,
      PCOUT(13) => blk00000001_sig000008ff,
      PCOUT(12) => blk00000001_sig000008fe,
      PCOUT(11) => blk00000001_sig000008fd,
      PCOUT(10) => blk00000001_sig000008fc,
      PCOUT(9) => blk00000001_sig000008fb,
      PCOUT(8) => blk00000001_sig000008fa,
      PCOUT(7) => blk00000001_sig000008f9,
      PCOUT(6) => blk00000001_sig000008f8,
      PCOUT(5) => blk00000001_sig000008f7,
      PCOUT(4) => blk00000001_sig000008f6,
      PCOUT(3) => blk00000001_sig000008f5,
      PCOUT(2) => blk00000001_sig000008f4,
      PCOUT(1) => blk00000001_sig000008f3,
      PCOUT(0) => blk00000001_sig000008f2,
      ACOUT(29) => NLW_blk00000001_blk00000d4a_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d4a_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d4a_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d4a_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d4a_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d4a_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d4a_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d4a_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d4a_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d4a_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d4a_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d4a_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d4a_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d4a_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d4a_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d4a_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d4a_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d4a_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d4a_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d4a_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d4a_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d4a_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d4a_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d4a_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d4a_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d4a_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d4a_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d4a_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d4a_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d4a_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d4a_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d4a_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d4a_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d4a_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d4a_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d4a_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d4a_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d4a_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d4a_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d4a_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d4a_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d4a_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d4a_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d4a_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d4a_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d4a_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d4a_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d4a_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d4a_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d4a_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d4a_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d4a_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d4a_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d4a_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d4a_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d4a_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d4a_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d4a_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d4a_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d4a_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d4a_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d4a_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d4a_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d4a_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d4a_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d4a_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d4a_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d4a_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d4a_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d4a_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d4a_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d4a_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d4a_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d4a_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d4a_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d4a_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d4a_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d4a_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d4a_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d4a_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d4a_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d4a_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d4a_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d4a_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d4a_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d4a_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d4a_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d4a_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d4a_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d4a_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d4a_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d4a_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d4a_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d4a_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d4a_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d4a_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d4a_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d4a_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d4a_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d4a_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d49 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d49_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d49_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d49_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d49_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d49_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d49_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig00000921,
      PCIN(46) => blk00000001_sig00000920,
      PCIN(45) => blk00000001_sig0000091f,
      PCIN(44) => blk00000001_sig0000091e,
      PCIN(43) => blk00000001_sig0000091d,
      PCIN(42) => blk00000001_sig0000091c,
      PCIN(41) => blk00000001_sig0000091b,
      PCIN(40) => blk00000001_sig0000091a,
      PCIN(39) => blk00000001_sig00000919,
      PCIN(38) => blk00000001_sig00000918,
      PCIN(37) => blk00000001_sig00000917,
      PCIN(36) => blk00000001_sig00000916,
      PCIN(35) => blk00000001_sig00000915,
      PCIN(34) => blk00000001_sig00000914,
      PCIN(33) => blk00000001_sig00000913,
      PCIN(32) => blk00000001_sig00000912,
      PCIN(31) => blk00000001_sig00000911,
      PCIN(30) => blk00000001_sig00000910,
      PCIN(29) => blk00000001_sig0000090f,
      PCIN(28) => blk00000001_sig0000090e,
      PCIN(27) => blk00000001_sig0000090d,
      PCIN(26) => blk00000001_sig0000090c,
      PCIN(25) => blk00000001_sig0000090b,
      PCIN(24) => blk00000001_sig0000090a,
      PCIN(23) => blk00000001_sig00000909,
      PCIN(22) => blk00000001_sig00000908,
      PCIN(21) => blk00000001_sig00000907,
      PCIN(20) => blk00000001_sig00000906,
      PCIN(19) => blk00000001_sig00000905,
      PCIN(18) => blk00000001_sig00000904,
      PCIN(17) => blk00000001_sig00000903,
      PCIN(16) => blk00000001_sig00000902,
      PCIN(15) => blk00000001_sig00000901,
      PCIN(14) => blk00000001_sig00000900,
      PCIN(13) => blk00000001_sig000008ff,
      PCIN(12) => blk00000001_sig000008fe,
      PCIN(11) => blk00000001_sig000008fd,
      PCIN(10) => blk00000001_sig000008fc,
      PCIN(9) => blk00000001_sig000008fb,
      PCIN(8) => blk00000001_sig000008fa,
      PCIN(7) => blk00000001_sig000008f9,
      PCIN(6) => blk00000001_sig000008f8,
      PCIN(5) => blk00000001_sig000008f7,
      PCIN(4) => blk00000001_sig000008f6,
      PCIN(3) => blk00000001_sig000008f5,
      PCIN(2) => blk00000001_sig000008f4,
      PCIN(1) => blk00000001_sig000008f3,
      PCIN(0) => blk00000001_sig000008f2,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig000007d7,
      B(16) => blk00000001_sig000007d7,
      B(15) => blk00000001_sig000007d7,
      B(14) => blk00000001_sig000007d6,
      B(13) => blk00000001_sig000007d5,
      B(12) => blk00000001_sig000007d4,
      B(11) => blk00000001_sig000007d3,
      B(10) => blk00000001_sig000007d2,
      B(9) => blk00000001_sig000007d1,
      B(8) => blk00000001_sig000007d0,
      B(7) => blk00000001_sig000007cf,
      B(6) => blk00000001_sig000007ce,
      B(5) => blk00000001_sig000007cd,
      B(4) => blk00000001_sig000007cc,
      B(3) => blk00000001_sig000007cb,
      B(2) => blk00000001_sig000007ca,
      B(1) => blk00000001_sig000007c9,
      B(0) => blk00000001_sig000007c8,
      P(47) => NLW_blk00000001_blk00000d49_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d49_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d49_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d49_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d49_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d49_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d49_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d49_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d49_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d49_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d49_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d49_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d49_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d49_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d49_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d49_P_32_UNCONNECTED,
      P(31) => blk00000001_sig00000741,
      P(30) => blk00000001_sig00000740,
      P(29) => blk00000001_sig0000073f,
      P(28) => blk00000001_sig0000073e,
      P(27) => blk00000001_sig0000073d,
      P(26) => blk00000001_sig0000073c,
      P(25) => blk00000001_sig0000073b,
      P(24) => blk00000001_sig0000073a,
      P(23) => blk00000001_sig00000739,
      P(22) => blk00000001_sig00000738,
      P(21) => blk00000001_sig00000737,
      P(20) => blk00000001_sig00000736,
      P(19) => blk00000001_sig00000735,
      P(18) => blk00000001_sig00000734,
      P(17) => blk00000001_sig00000733,
      P(16) => blk00000001_sig00000732,
      P(15) => blk00000001_sig00000731,
      P(14) => blk00000001_sig00000730,
      P(13) => blk00000001_sig0000072f,
      P(12) => blk00000001_sig0000072e,
      P(11) => NLW_blk00000001_blk00000d49_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d49_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d49_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d49_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d49_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d49_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d49_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d49_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d49_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d49_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d49_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d49_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig00000809,
      A(23) => blk00000001_sig00000809,
      A(22) => blk00000001_sig00000809,
      A(21) => blk00000001_sig00000809,
      A(20) => blk00000001_sig00000809,
      A(19) => blk00000001_sig00000809,
      A(18) => blk00000001_sig00000809,
      A(17) => blk00000001_sig00000809,
      A(16) => blk00000001_sig00000809,
      A(15) => blk00000001_sig00000808,
      A(14) => blk00000001_sig00000807,
      A(13) => blk00000001_sig00000806,
      A(12) => blk00000001_sig00000805,
      A(11) => blk00000001_sig00000804,
      A(10) => blk00000001_sig00000803,
      A(9) => blk00000001_sig00000802,
      A(8) => blk00000001_sig00000801,
      A(7) => blk00000001_sig00000800,
      A(6) => blk00000001_sig000007ff,
      A(5) => blk00000001_sig000007fe,
      A(4) => blk00000001_sig000007fd,
      A(3) => blk00000001_sig000007fc,
      A(2) => blk00000001_sig000007fb,
      A(1) => blk00000001_sig000007fa,
      A(0) => blk00000001_sig000007f9,
      PCOUT(47) => NLW_blk00000001_blk00000d49_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d49_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d49_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d49_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d49_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d49_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d49_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d49_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d49_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d49_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d49_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d49_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d49_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d49_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d49_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d49_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d49_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d49_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d49_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d49_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d49_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d49_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d49_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d49_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d49_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d49_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d49_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d49_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d49_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d49_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d49_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d49_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d49_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d49_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d49_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d49_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d49_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d49_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d49_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d49_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d49_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d49_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d49_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d49_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d49_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d49_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d49_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d49_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d49_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d49_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d49_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d49_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d49_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d49_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d49_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d49_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d49_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d49_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d49_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d49_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d49_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d49_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d49_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d49_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d49_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d49_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d49_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d49_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d49_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d49_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d49_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d49_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d49_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d49_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d49_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d49_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d49_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d49_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d49_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d49_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d49_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d49_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d49_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d49_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d49_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d49_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d49_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d49_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d49_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d49_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d49_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d49_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d49_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d49_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d49_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d49_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d49_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d49_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d49_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d49_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d48 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d48_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d48_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d48_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d48_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d48_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d48_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig000008af,
      ALUMODE(0) => blk00000001_sig000008af,
      B(17) => blk00000001_sig000008cf,
      B(16) => blk00000001_sig000008cf,
      B(15) => blk00000001_sig000008cf,
      B(14) => blk00000001_sig000008ce,
      B(13) => blk00000001_sig000008cd,
      B(12) => blk00000001_sig000008cc,
      B(11) => blk00000001_sig000008cb,
      B(10) => blk00000001_sig000008ca,
      B(9) => blk00000001_sig000008c9,
      B(8) => blk00000001_sig000008c8,
      B(7) => blk00000001_sig000008c7,
      B(6) => blk00000001_sig000008c6,
      B(5) => blk00000001_sig000008c5,
      B(4) => blk00000001_sig000008c4,
      B(3) => blk00000001_sig000008c3,
      B(2) => blk00000001_sig000008c2,
      B(1) => blk00000001_sig000008c1,
      B(0) => blk00000001_sig000008c0,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000008f1,
      A(23) => blk00000001_sig000008f1,
      A(22) => blk00000001_sig000008f1,
      A(21) => blk00000001_sig000008f1,
      A(20) => blk00000001_sig000008f1,
      A(19) => blk00000001_sig000008f1,
      A(18) => blk00000001_sig000008f1,
      A(17) => blk00000001_sig000008f1,
      A(16) => blk00000001_sig000008f1,
      A(15) => blk00000001_sig000008f0,
      A(14) => blk00000001_sig000008ef,
      A(13) => blk00000001_sig000008ee,
      A(12) => blk00000001_sig000008ed,
      A(11) => blk00000001_sig000008ec,
      A(10) => blk00000001_sig000008eb,
      A(9) => blk00000001_sig000008ea,
      A(8) => blk00000001_sig000008e9,
      A(7) => blk00000001_sig000008e8,
      A(6) => blk00000001_sig000008e7,
      A(5) => blk00000001_sig000008e6,
      A(4) => blk00000001_sig000008e5,
      A(3) => blk00000001_sig000008e4,
      A(2) => blk00000001_sig000008e3,
      A(1) => blk00000001_sig000008e2,
      A(0) => blk00000001_sig000008e1,
      PCOUT(47) => blk00000001_sig000008ad,
      PCOUT(46) => blk00000001_sig000008ac,
      PCOUT(45) => blk00000001_sig000008ab,
      PCOUT(44) => blk00000001_sig000008aa,
      PCOUT(43) => blk00000001_sig000008a9,
      PCOUT(42) => blk00000001_sig000008a8,
      PCOUT(41) => blk00000001_sig000008a7,
      PCOUT(40) => blk00000001_sig000008a6,
      PCOUT(39) => blk00000001_sig000008a5,
      PCOUT(38) => blk00000001_sig000008a4,
      PCOUT(37) => blk00000001_sig000008a3,
      PCOUT(36) => blk00000001_sig000008a2,
      PCOUT(35) => blk00000001_sig000008a1,
      PCOUT(34) => blk00000001_sig000008a0,
      PCOUT(33) => blk00000001_sig0000089f,
      PCOUT(32) => blk00000001_sig0000089e,
      PCOUT(31) => blk00000001_sig0000089d,
      PCOUT(30) => blk00000001_sig0000089c,
      PCOUT(29) => blk00000001_sig0000089b,
      PCOUT(28) => blk00000001_sig0000089a,
      PCOUT(27) => blk00000001_sig00000899,
      PCOUT(26) => blk00000001_sig00000898,
      PCOUT(25) => blk00000001_sig00000897,
      PCOUT(24) => blk00000001_sig00000896,
      PCOUT(23) => blk00000001_sig00000895,
      PCOUT(22) => blk00000001_sig00000894,
      PCOUT(21) => blk00000001_sig00000893,
      PCOUT(20) => blk00000001_sig00000892,
      PCOUT(19) => blk00000001_sig00000891,
      PCOUT(18) => blk00000001_sig00000890,
      PCOUT(17) => blk00000001_sig0000088f,
      PCOUT(16) => blk00000001_sig0000088e,
      PCOUT(15) => blk00000001_sig0000088d,
      PCOUT(14) => blk00000001_sig0000088c,
      PCOUT(13) => blk00000001_sig0000088b,
      PCOUT(12) => blk00000001_sig0000088a,
      PCOUT(11) => blk00000001_sig00000889,
      PCOUT(10) => blk00000001_sig00000888,
      PCOUT(9) => blk00000001_sig00000887,
      PCOUT(8) => blk00000001_sig00000886,
      PCOUT(7) => blk00000001_sig00000885,
      PCOUT(6) => blk00000001_sig00000884,
      PCOUT(5) => blk00000001_sig00000883,
      PCOUT(4) => blk00000001_sig00000882,
      PCOUT(3) => blk00000001_sig00000881,
      PCOUT(2) => blk00000001_sig00000880,
      PCOUT(1) => blk00000001_sig0000087f,
      PCOUT(0) => blk00000001_sig0000087e,
      ACOUT(29) => NLW_blk00000001_blk00000d48_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d48_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d48_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d48_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d48_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d48_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d48_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d48_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d48_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d48_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d48_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d48_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d48_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d48_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d48_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d48_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d48_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d48_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d48_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d48_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d48_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d48_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d48_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d48_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d48_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d48_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d48_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d48_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d48_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d48_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d48_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d48_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d48_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d48_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d48_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d48_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d48_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d48_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d48_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d48_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d48_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d48_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d48_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d48_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d48_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d48_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d48_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d48_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d48_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d48_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d48_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d48_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d48_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d48_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d48_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d48_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d48_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d48_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d48_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d48_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d48_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d48_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d48_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d48_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d48_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d48_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d48_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d48_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d48_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d48_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d48_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d48_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d48_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d48_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d48_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d48_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d48_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d48_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d48_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d48_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d48_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d48_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d48_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d48_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d48_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d48_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d48_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d48_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d48_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d48_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d48_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d48_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d48_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d48_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d48_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d48_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d48_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d48_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d48_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d48_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d47 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d47_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d47_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d47_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d47_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d47_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d47_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig000008ad,
      PCIN(46) => blk00000001_sig000008ac,
      PCIN(45) => blk00000001_sig000008ab,
      PCIN(44) => blk00000001_sig000008aa,
      PCIN(43) => blk00000001_sig000008a9,
      PCIN(42) => blk00000001_sig000008a8,
      PCIN(41) => blk00000001_sig000008a7,
      PCIN(40) => blk00000001_sig000008a6,
      PCIN(39) => blk00000001_sig000008a5,
      PCIN(38) => blk00000001_sig000008a4,
      PCIN(37) => blk00000001_sig000008a3,
      PCIN(36) => blk00000001_sig000008a2,
      PCIN(35) => blk00000001_sig000008a1,
      PCIN(34) => blk00000001_sig000008a0,
      PCIN(33) => blk00000001_sig0000089f,
      PCIN(32) => blk00000001_sig0000089e,
      PCIN(31) => blk00000001_sig0000089d,
      PCIN(30) => blk00000001_sig0000089c,
      PCIN(29) => blk00000001_sig0000089b,
      PCIN(28) => blk00000001_sig0000089a,
      PCIN(27) => blk00000001_sig00000899,
      PCIN(26) => blk00000001_sig00000898,
      PCIN(25) => blk00000001_sig00000897,
      PCIN(24) => blk00000001_sig00000896,
      PCIN(23) => blk00000001_sig00000895,
      PCIN(22) => blk00000001_sig00000894,
      PCIN(21) => blk00000001_sig00000893,
      PCIN(20) => blk00000001_sig00000892,
      PCIN(19) => blk00000001_sig00000891,
      PCIN(18) => blk00000001_sig00000890,
      PCIN(17) => blk00000001_sig0000088f,
      PCIN(16) => blk00000001_sig0000088e,
      PCIN(15) => blk00000001_sig0000088d,
      PCIN(14) => blk00000001_sig0000088c,
      PCIN(13) => blk00000001_sig0000088b,
      PCIN(12) => blk00000001_sig0000088a,
      PCIN(11) => blk00000001_sig00000889,
      PCIN(10) => blk00000001_sig00000888,
      PCIN(9) => blk00000001_sig00000887,
      PCIN(8) => blk00000001_sig00000886,
      PCIN(7) => blk00000001_sig00000885,
      PCIN(6) => blk00000001_sig00000884,
      PCIN(5) => blk00000001_sig00000883,
      PCIN(4) => blk00000001_sig00000882,
      PCIN(3) => blk00000001_sig00000881,
      PCIN(2) => blk00000001_sig00000880,
      PCIN(1) => blk00000001_sig0000087f,
      PCIN(0) => blk00000001_sig0000087e,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig0000087d,
      ALUMODE(0) => blk00000001_sig0000087d,
      B(17) => blk00000001_sig000008bf,
      B(16) => blk00000001_sig000008bf,
      B(15) => blk00000001_sig000008bf,
      B(14) => blk00000001_sig000008be,
      B(13) => blk00000001_sig000008bd,
      B(12) => blk00000001_sig000008bc,
      B(11) => blk00000001_sig000008bb,
      B(10) => blk00000001_sig000008ba,
      B(9) => blk00000001_sig000008b9,
      B(8) => blk00000001_sig000008b8,
      B(7) => blk00000001_sig000008b7,
      B(6) => blk00000001_sig000008b6,
      B(5) => blk00000001_sig000008b5,
      B(4) => blk00000001_sig000008b4,
      B(3) => blk00000001_sig000008b3,
      B(2) => blk00000001_sig000008b2,
      B(1) => blk00000001_sig000008b1,
      B(0) => blk00000001_sig000008b0,
      P(47) => NLW_blk00000001_blk00000d47_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d47_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d47_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d47_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d47_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d47_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d47_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d47_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d47_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d47_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d47_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d47_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d47_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d47_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d47_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d47_P_32_UNCONNECTED,
      P(31) => blk00000001_sig00000705,
      P(30) => blk00000001_sig00000704,
      P(29) => blk00000001_sig00000703,
      P(28) => blk00000001_sig00000702,
      P(27) => blk00000001_sig00000701,
      P(26) => blk00000001_sig00000700,
      P(25) => blk00000001_sig000006ff,
      P(24) => blk00000001_sig000006fe,
      P(23) => blk00000001_sig000006fd,
      P(22) => blk00000001_sig000006fc,
      P(21) => blk00000001_sig000006fb,
      P(20) => blk00000001_sig000006fa,
      P(19) => blk00000001_sig000006f9,
      P(18) => blk00000001_sig000006f8,
      P(17) => blk00000001_sig000006f7,
      P(16) => blk00000001_sig000006f6,
      P(15) => blk00000001_sig000006f5,
      P(14) => blk00000001_sig000006f4,
      P(13) => blk00000001_sig000006f3,
      P(12) => blk00000001_sig000006f2,
      P(11) => NLW_blk00000001_blk00000d47_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d47_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d47_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d47_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d47_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d47_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d47_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d47_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d47_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d47_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d47_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d47_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000008e0,
      A(23) => blk00000001_sig000008e0,
      A(22) => blk00000001_sig000008e0,
      A(21) => blk00000001_sig000008e0,
      A(20) => blk00000001_sig000008e0,
      A(19) => blk00000001_sig000008e0,
      A(18) => blk00000001_sig000008e0,
      A(17) => blk00000001_sig000008e0,
      A(16) => blk00000001_sig000008e0,
      A(15) => blk00000001_sig000008df,
      A(14) => blk00000001_sig000008de,
      A(13) => blk00000001_sig000008dd,
      A(12) => blk00000001_sig000008dc,
      A(11) => blk00000001_sig000008db,
      A(10) => blk00000001_sig000008da,
      A(9) => blk00000001_sig000008d9,
      A(8) => blk00000001_sig000008d8,
      A(7) => blk00000001_sig000008d7,
      A(6) => blk00000001_sig000008d6,
      A(5) => blk00000001_sig000008d5,
      A(4) => blk00000001_sig000008d4,
      A(3) => blk00000001_sig000008d3,
      A(2) => blk00000001_sig000008d2,
      A(1) => blk00000001_sig000008d1,
      A(0) => blk00000001_sig000008d0,
      PCOUT(47) => NLW_blk00000001_blk00000d47_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d47_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d47_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d47_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d47_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d47_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d47_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d47_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d47_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d47_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d47_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d47_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d47_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d47_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d47_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d47_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d47_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d47_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d47_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d47_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d47_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d47_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d47_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d47_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d47_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d47_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d47_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d47_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d47_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d47_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d47_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d47_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d47_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d47_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d47_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d47_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d47_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d47_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d47_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d47_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d47_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d47_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d47_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d47_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d47_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d47_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d47_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d47_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d47_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d47_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d47_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d47_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d47_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d47_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d47_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d47_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d47_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d47_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d47_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d47_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d47_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d47_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d47_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d47_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d47_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d47_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d47_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d47_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d47_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d47_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d47_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d47_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d47_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d47_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d47_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d47_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d47_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d47_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d47_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d47_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d47_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d47_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d47_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d47_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d47_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d47_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d47_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d47_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d47_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d47_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d47_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d47_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d47_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d47_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d47_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d47_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d47_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d47_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d47_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d47_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d46 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d46_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d46_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d46_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d46_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d46_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d46_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig0000085a,
      B(16) => blk00000001_sig0000085a,
      B(15) => blk00000001_sig0000085a,
      B(14) => blk00000001_sig00000859,
      B(13) => blk00000001_sig00000858,
      B(12) => blk00000001_sig00000857,
      B(11) => blk00000001_sig00000856,
      B(10) => blk00000001_sig00000855,
      B(9) => blk00000001_sig00000854,
      B(8) => blk00000001_sig00000853,
      B(7) => blk00000001_sig00000852,
      B(6) => blk00000001_sig00000851,
      B(5) => blk00000001_sig00000850,
      B(4) => blk00000001_sig0000084f,
      B(3) => blk00000001_sig0000084e,
      B(2) => blk00000001_sig0000084d,
      B(1) => blk00000001_sig0000084c,
      B(0) => blk00000001_sig0000084b,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig0000087c,
      A(23) => blk00000001_sig0000087c,
      A(22) => blk00000001_sig0000087c,
      A(21) => blk00000001_sig0000087c,
      A(20) => blk00000001_sig0000087c,
      A(19) => blk00000001_sig0000087c,
      A(18) => blk00000001_sig0000087c,
      A(17) => blk00000001_sig0000087c,
      A(16) => blk00000001_sig0000087c,
      A(15) => blk00000001_sig0000087b,
      A(14) => blk00000001_sig0000087a,
      A(13) => blk00000001_sig00000879,
      A(12) => blk00000001_sig00000878,
      A(11) => blk00000001_sig00000877,
      A(10) => blk00000001_sig00000876,
      A(9) => blk00000001_sig00000875,
      A(8) => blk00000001_sig00000874,
      A(7) => blk00000001_sig00000873,
      A(6) => blk00000001_sig00000872,
      A(5) => blk00000001_sig00000871,
      A(4) => blk00000001_sig00000870,
      A(3) => blk00000001_sig0000086f,
      A(2) => blk00000001_sig0000086e,
      A(1) => blk00000001_sig0000086d,
      A(0) => blk00000001_sig0000086c,
      PCOUT(47) => blk00000001_sig0000083a,
      PCOUT(46) => blk00000001_sig00000839,
      PCOUT(45) => blk00000001_sig00000838,
      PCOUT(44) => blk00000001_sig00000837,
      PCOUT(43) => blk00000001_sig00000836,
      PCOUT(42) => blk00000001_sig00000835,
      PCOUT(41) => blk00000001_sig00000834,
      PCOUT(40) => blk00000001_sig00000833,
      PCOUT(39) => blk00000001_sig00000832,
      PCOUT(38) => blk00000001_sig00000831,
      PCOUT(37) => blk00000001_sig00000830,
      PCOUT(36) => blk00000001_sig0000082f,
      PCOUT(35) => blk00000001_sig0000082e,
      PCOUT(34) => blk00000001_sig0000082d,
      PCOUT(33) => blk00000001_sig0000082c,
      PCOUT(32) => blk00000001_sig0000082b,
      PCOUT(31) => blk00000001_sig0000082a,
      PCOUT(30) => blk00000001_sig00000829,
      PCOUT(29) => blk00000001_sig00000828,
      PCOUT(28) => blk00000001_sig00000827,
      PCOUT(27) => blk00000001_sig00000826,
      PCOUT(26) => blk00000001_sig00000825,
      PCOUT(25) => blk00000001_sig00000824,
      PCOUT(24) => blk00000001_sig00000823,
      PCOUT(23) => blk00000001_sig00000822,
      PCOUT(22) => blk00000001_sig00000821,
      PCOUT(21) => blk00000001_sig00000820,
      PCOUT(20) => blk00000001_sig0000081f,
      PCOUT(19) => blk00000001_sig0000081e,
      PCOUT(18) => blk00000001_sig0000081d,
      PCOUT(17) => blk00000001_sig0000081c,
      PCOUT(16) => blk00000001_sig0000081b,
      PCOUT(15) => blk00000001_sig0000081a,
      PCOUT(14) => blk00000001_sig00000819,
      PCOUT(13) => blk00000001_sig00000818,
      PCOUT(12) => blk00000001_sig00000817,
      PCOUT(11) => blk00000001_sig00000816,
      PCOUT(10) => blk00000001_sig00000815,
      PCOUT(9) => blk00000001_sig00000814,
      PCOUT(8) => blk00000001_sig00000813,
      PCOUT(7) => blk00000001_sig00000812,
      PCOUT(6) => blk00000001_sig00000811,
      PCOUT(5) => blk00000001_sig00000810,
      PCOUT(4) => blk00000001_sig0000080f,
      PCOUT(3) => blk00000001_sig0000080e,
      PCOUT(2) => blk00000001_sig0000080d,
      PCOUT(1) => blk00000001_sig0000080c,
      PCOUT(0) => blk00000001_sig0000080b,
      ACOUT(29) => NLW_blk00000001_blk00000d46_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d46_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d46_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d46_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d46_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d46_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d46_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d46_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d46_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d46_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d46_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d46_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d46_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d46_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d46_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d46_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d46_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d46_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d46_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d46_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d46_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d46_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d46_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d46_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d46_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d46_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d46_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d46_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d46_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d46_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d46_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d46_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d46_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d46_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d46_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d46_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d46_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d46_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d46_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d46_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d46_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d46_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d46_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d46_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d46_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d46_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d46_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d46_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d46_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d46_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d46_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d46_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d46_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d46_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d46_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d46_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d46_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d46_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d46_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d46_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d46_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d46_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d46_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d46_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d46_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d46_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d46_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d46_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d46_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d46_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d46_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d46_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d46_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d46_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d46_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d46_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d46_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d46_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d46_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d46_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d46_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d46_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d46_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d46_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d46_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d46_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d46_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d46_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d46_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d46_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d46_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d46_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d46_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d46_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d46_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d46_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d46_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d46_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d46_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d46_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d45 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d45_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d45_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d45_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d45_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d45_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d45_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig0000083a,
      PCIN(46) => blk00000001_sig00000839,
      PCIN(45) => blk00000001_sig00000838,
      PCIN(44) => blk00000001_sig00000837,
      PCIN(43) => blk00000001_sig00000836,
      PCIN(42) => blk00000001_sig00000835,
      PCIN(41) => blk00000001_sig00000834,
      PCIN(40) => blk00000001_sig00000833,
      PCIN(39) => blk00000001_sig00000832,
      PCIN(38) => blk00000001_sig00000831,
      PCIN(37) => blk00000001_sig00000830,
      PCIN(36) => blk00000001_sig0000082f,
      PCIN(35) => blk00000001_sig0000082e,
      PCIN(34) => blk00000001_sig0000082d,
      PCIN(33) => blk00000001_sig0000082c,
      PCIN(32) => blk00000001_sig0000082b,
      PCIN(31) => blk00000001_sig0000082a,
      PCIN(30) => blk00000001_sig00000829,
      PCIN(29) => blk00000001_sig00000828,
      PCIN(28) => blk00000001_sig00000827,
      PCIN(27) => blk00000001_sig00000826,
      PCIN(26) => blk00000001_sig00000825,
      PCIN(25) => blk00000001_sig00000824,
      PCIN(24) => blk00000001_sig00000823,
      PCIN(23) => blk00000001_sig00000822,
      PCIN(22) => blk00000001_sig00000821,
      PCIN(21) => blk00000001_sig00000820,
      PCIN(20) => blk00000001_sig0000081f,
      PCIN(19) => blk00000001_sig0000081e,
      PCIN(18) => blk00000001_sig0000081d,
      PCIN(17) => blk00000001_sig0000081c,
      PCIN(16) => blk00000001_sig0000081b,
      PCIN(15) => blk00000001_sig0000081a,
      PCIN(14) => blk00000001_sig00000819,
      PCIN(13) => blk00000001_sig00000818,
      PCIN(12) => blk00000001_sig00000817,
      PCIN(11) => blk00000001_sig00000816,
      PCIN(10) => blk00000001_sig00000815,
      PCIN(9) => blk00000001_sig00000814,
      PCIN(8) => blk00000001_sig00000813,
      PCIN(7) => blk00000001_sig00000812,
      PCIN(6) => blk00000001_sig00000811,
      PCIN(5) => blk00000001_sig00000810,
      PCIN(4) => blk00000001_sig0000080f,
      PCIN(3) => blk00000001_sig0000080e,
      PCIN(2) => blk00000001_sig0000080d,
      PCIN(1) => blk00000001_sig0000080c,
      PCIN(0) => blk00000001_sig0000080b,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig0000080a,
      ALUMODE(0) => blk00000001_sig0000080a,
      B(17) => blk00000001_sig0000084a,
      B(16) => blk00000001_sig0000084a,
      B(15) => blk00000001_sig0000084a,
      B(14) => blk00000001_sig00000849,
      B(13) => blk00000001_sig00000848,
      B(12) => blk00000001_sig00000847,
      B(11) => blk00000001_sig00000846,
      B(10) => blk00000001_sig00000845,
      B(9) => blk00000001_sig00000844,
      B(8) => blk00000001_sig00000843,
      B(7) => blk00000001_sig00000842,
      B(6) => blk00000001_sig00000841,
      B(5) => blk00000001_sig00000840,
      B(4) => blk00000001_sig0000083f,
      B(3) => blk00000001_sig0000083e,
      B(2) => blk00000001_sig0000083d,
      B(1) => blk00000001_sig0000083c,
      B(0) => blk00000001_sig0000083b,
      P(47) => NLW_blk00000001_blk00000d45_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d45_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d45_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d45_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d45_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d45_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d45_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d45_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d45_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d45_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d45_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d45_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d45_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d45_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d45_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d45_P_32_UNCONNECTED,
      P(31) => blk00000001_sig0000072d,
      P(30) => blk00000001_sig0000072c,
      P(29) => blk00000001_sig0000072b,
      P(28) => blk00000001_sig0000072a,
      P(27) => blk00000001_sig00000729,
      P(26) => blk00000001_sig00000728,
      P(25) => blk00000001_sig00000727,
      P(24) => blk00000001_sig00000726,
      P(23) => blk00000001_sig00000725,
      P(22) => blk00000001_sig00000724,
      P(21) => blk00000001_sig00000723,
      P(20) => blk00000001_sig00000722,
      P(19) => blk00000001_sig00000721,
      P(18) => blk00000001_sig00000720,
      P(17) => blk00000001_sig0000071f,
      P(16) => blk00000001_sig0000071e,
      P(15) => blk00000001_sig0000071d,
      P(14) => blk00000001_sig0000071c,
      P(13) => blk00000001_sig0000071b,
      P(12) => blk00000001_sig0000071a,
      P(11) => NLW_blk00000001_blk00000d45_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d45_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d45_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d45_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d45_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d45_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d45_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d45_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d45_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d45_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d45_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d45_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig0000086b,
      A(23) => blk00000001_sig0000086b,
      A(22) => blk00000001_sig0000086b,
      A(21) => blk00000001_sig0000086b,
      A(20) => blk00000001_sig0000086b,
      A(19) => blk00000001_sig0000086b,
      A(18) => blk00000001_sig0000086b,
      A(17) => blk00000001_sig0000086b,
      A(16) => blk00000001_sig0000086b,
      A(15) => blk00000001_sig0000086a,
      A(14) => blk00000001_sig00000869,
      A(13) => blk00000001_sig00000868,
      A(12) => blk00000001_sig00000867,
      A(11) => blk00000001_sig00000866,
      A(10) => blk00000001_sig00000865,
      A(9) => blk00000001_sig00000864,
      A(8) => blk00000001_sig00000863,
      A(7) => blk00000001_sig00000862,
      A(6) => blk00000001_sig00000861,
      A(5) => blk00000001_sig00000860,
      A(4) => blk00000001_sig0000085f,
      A(3) => blk00000001_sig0000085e,
      A(2) => blk00000001_sig0000085d,
      A(1) => blk00000001_sig0000085c,
      A(0) => blk00000001_sig0000085b,
      PCOUT(47) => NLW_blk00000001_blk00000d45_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d45_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d45_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d45_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d45_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d45_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d45_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d45_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d45_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d45_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d45_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d45_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d45_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d45_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d45_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d45_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d45_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d45_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d45_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d45_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d45_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d45_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d45_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d45_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d45_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d45_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d45_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d45_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d45_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d45_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d45_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d45_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d45_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d45_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d45_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d45_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d45_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d45_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d45_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d45_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d45_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d45_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d45_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d45_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d45_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d45_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d45_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d45_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d45_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d45_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d45_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d45_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d45_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d45_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d45_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d45_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d45_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d45_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d45_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d45_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d45_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d45_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d45_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d45_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d45_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d45_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d45_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d45_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d45_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d45_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d45_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d45_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d45_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d45_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d45_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d45_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d45_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d45_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d45_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d45_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d45_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d45_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d45_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d45_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d45_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d45_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d45_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d45_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d45_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d45_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d45_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d45_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d45_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d45_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d45_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d45_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d45_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d45_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d45_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d45_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d44 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d44_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNOUT => NLW_blk00000001_blk00000d44_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d44_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d44_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d44_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d44_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      B(17) => blk00000001_sig000007e7,
      B(16) => blk00000001_sig000007e7,
      B(15) => blk00000001_sig000007e7,
      B(14) => blk00000001_sig000007e6,
      B(13) => blk00000001_sig000007e5,
      B(12) => blk00000001_sig000007e4,
      B(11) => blk00000001_sig000007e3,
      B(10) => blk00000001_sig000007e2,
      B(9) => blk00000001_sig000007e1,
      B(8) => blk00000001_sig000007e0,
      B(7) => blk00000001_sig000007df,
      B(6) => blk00000001_sig000007de,
      B(5) => blk00000001_sig000007dd,
      B(4) => blk00000001_sig000007dc,
      B(3) => blk00000001_sig000007db,
      B(2) => blk00000001_sig000007da,
      B(1) => blk00000001_sig000007d9,
      B(0) => blk00000001_sig000007d8,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig00000809,
      A(23) => blk00000001_sig00000809,
      A(22) => blk00000001_sig00000809,
      A(21) => blk00000001_sig00000809,
      A(20) => blk00000001_sig00000809,
      A(19) => blk00000001_sig00000809,
      A(18) => blk00000001_sig00000809,
      A(17) => blk00000001_sig00000809,
      A(16) => blk00000001_sig00000809,
      A(15) => blk00000001_sig00000808,
      A(14) => blk00000001_sig00000807,
      A(13) => blk00000001_sig00000806,
      A(12) => blk00000001_sig00000805,
      A(11) => blk00000001_sig00000804,
      A(10) => blk00000001_sig00000803,
      A(9) => blk00000001_sig00000802,
      A(8) => blk00000001_sig00000801,
      A(7) => blk00000001_sig00000800,
      A(6) => blk00000001_sig000007ff,
      A(5) => blk00000001_sig000007fe,
      A(4) => blk00000001_sig000007fd,
      A(3) => blk00000001_sig000007fc,
      A(2) => blk00000001_sig000007fb,
      A(1) => blk00000001_sig000007fa,
      A(0) => blk00000001_sig000007f9,
      PCOUT(47) => blk00000001_sig000007c6,
      PCOUT(46) => blk00000001_sig000007c5,
      PCOUT(45) => blk00000001_sig000007c4,
      PCOUT(44) => blk00000001_sig000007c3,
      PCOUT(43) => blk00000001_sig000007c2,
      PCOUT(42) => blk00000001_sig000007c1,
      PCOUT(41) => blk00000001_sig000007c0,
      PCOUT(40) => blk00000001_sig000007bf,
      PCOUT(39) => blk00000001_sig000007be,
      PCOUT(38) => blk00000001_sig000007bd,
      PCOUT(37) => blk00000001_sig000007bc,
      PCOUT(36) => blk00000001_sig000007bb,
      PCOUT(35) => blk00000001_sig000007ba,
      PCOUT(34) => blk00000001_sig000007b9,
      PCOUT(33) => blk00000001_sig000007b8,
      PCOUT(32) => blk00000001_sig000007b7,
      PCOUT(31) => blk00000001_sig000007b6,
      PCOUT(30) => blk00000001_sig000007b5,
      PCOUT(29) => blk00000001_sig000007b4,
      PCOUT(28) => blk00000001_sig000007b3,
      PCOUT(27) => blk00000001_sig000007b2,
      PCOUT(26) => blk00000001_sig000007b1,
      PCOUT(25) => blk00000001_sig000007b0,
      PCOUT(24) => blk00000001_sig000007af,
      PCOUT(23) => blk00000001_sig000007ae,
      PCOUT(22) => blk00000001_sig000007ad,
      PCOUT(21) => blk00000001_sig000007ac,
      PCOUT(20) => blk00000001_sig000007ab,
      PCOUT(19) => blk00000001_sig000007aa,
      PCOUT(18) => blk00000001_sig000007a9,
      PCOUT(17) => blk00000001_sig000007a8,
      PCOUT(16) => blk00000001_sig000007a7,
      PCOUT(15) => blk00000001_sig000007a6,
      PCOUT(14) => blk00000001_sig000007a5,
      PCOUT(13) => blk00000001_sig000007a4,
      PCOUT(12) => blk00000001_sig000007a3,
      PCOUT(11) => blk00000001_sig000007a2,
      PCOUT(10) => blk00000001_sig000007a1,
      PCOUT(9) => blk00000001_sig000007a0,
      PCOUT(8) => blk00000001_sig0000079f,
      PCOUT(7) => blk00000001_sig0000079e,
      PCOUT(6) => blk00000001_sig0000079d,
      PCOUT(5) => blk00000001_sig0000079c,
      PCOUT(4) => blk00000001_sig0000079b,
      PCOUT(3) => blk00000001_sig0000079a,
      PCOUT(2) => blk00000001_sig00000799,
      PCOUT(1) => blk00000001_sig00000798,
      PCOUT(0) => blk00000001_sig00000797,
      ACOUT(29) => NLW_blk00000001_blk00000d44_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d44_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d44_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d44_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d44_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d44_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d44_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d44_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d44_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d44_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d44_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d44_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d44_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d44_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d44_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d44_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d44_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d44_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d44_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d44_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d44_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d44_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d44_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d44_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d44_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d44_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d44_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d44_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d44_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d44_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => blk00000001_sig000000c0,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      PCIN(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      PCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYOUT(3) => NLW_blk00000001_blk00000d44_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d44_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d44_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d44_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d44_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d44_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d44_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d44_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d44_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d44_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d44_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d44_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d44_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d44_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d44_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d44_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d44_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d44_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d44_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d44_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d44_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d44_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk00000d44_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d44_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d44_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d44_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d44_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d44_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d44_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d44_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d44_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d44_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d44_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d44_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d44_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d44_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d44_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d44_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk00000d44_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk00000d44_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk00000d44_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk00000d44_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk00000d44_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk00000d44_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk00000d44_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk00000d44_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk00000d44_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk00000d44_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk00000d44_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk00000d44_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk00000d44_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk00000d44_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk00000d44_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk00000d44_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk00000d44_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk00000d44_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk00000d44_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk00000d44_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk00000d44_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d44_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d44_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d44_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d44_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d44_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d44_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d44_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d44_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d44_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d44_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d44_P_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d43 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000008e,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk00000d43_PATTERNBDETECT_UNCONNECTED,
      RSTC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB1 => blk00000001_sig0000008e,
      MULTSIGNOUT => NLW_blk00000001_blk00000d43_MULTSIGNOUT_UNCONNECTED,
      CEC => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      MULTSIGNIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEB2 => blk00000001_sig0000008e,
      RSTCTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEP => blk00000001_sig0000008e,
      CARRYCASCOUT => NLW_blk00000001_blk00000d43_CARRYCASCOUT_UNCONNECTED,
      RSTA => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CECARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      UNDERFLOW => NLW_blk00000001_blk00000d43_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk00000d43_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTALLCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEALUMODE => blk00000001_sig0000008e,
      CEA2 => blk00000001_sig0000008e,
      CEA1 => blk00000001_sig0000008e,
      RSTB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CEMULTCARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OVERFLOW => NLW_blk00000001_blk00000d43_OVERFLOW_UNCONNECTED,
      CECTRL => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYCASCIN => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTP => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CARRYINSEL(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(47) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(46) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(45) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(44) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(43) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(42) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(41) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(40) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(39) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(38) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(37) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(36) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(35) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(34) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(33) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(32) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(31) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(30) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      C(10) => blk00000001_sig000000c0,
      C(9) => blk00000001_sig000000c0,
      C(8) => blk00000001_sig000000c0,
      C(7) => blk00000001_sig000000c0,
      C(6) => blk00000001_sig000000c0,
      C(5) => blk00000001_sig000000c0,
      C(4) => blk00000001_sig000000c0,
      C(3) => blk00000001_sig000000c0,
      C(2) => blk00000001_sig000000c0,
      C(1) => blk00000001_sig000000c0,
      C(0) => blk00000001_sig000000c0,
      PCIN(47) => blk00000001_sig000007c6,
      PCIN(46) => blk00000001_sig000007c5,
      PCIN(45) => blk00000001_sig000007c4,
      PCIN(44) => blk00000001_sig000007c3,
      PCIN(43) => blk00000001_sig000007c2,
      PCIN(42) => blk00000001_sig000007c1,
      PCIN(41) => blk00000001_sig000007c0,
      PCIN(40) => blk00000001_sig000007bf,
      PCIN(39) => blk00000001_sig000007be,
      PCIN(38) => blk00000001_sig000007bd,
      PCIN(37) => blk00000001_sig000007bc,
      PCIN(36) => blk00000001_sig000007bb,
      PCIN(35) => blk00000001_sig000007ba,
      PCIN(34) => blk00000001_sig000007b9,
      PCIN(33) => blk00000001_sig000007b8,
      PCIN(32) => blk00000001_sig000007b7,
      PCIN(31) => blk00000001_sig000007b6,
      PCIN(30) => blk00000001_sig000007b5,
      PCIN(29) => blk00000001_sig000007b4,
      PCIN(28) => blk00000001_sig000007b3,
      PCIN(27) => blk00000001_sig000007b2,
      PCIN(26) => blk00000001_sig000007b1,
      PCIN(25) => blk00000001_sig000007b0,
      PCIN(24) => blk00000001_sig000007af,
      PCIN(23) => blk00000001_sig000007ae,
      PCIN(22) => blk00000001_sig000007ad,
      PCIN(21) => blk00000001_sig000007ac,
      PCIN(20) => blk00000001_sig000007ab,
      PCIN(19) => blk00000001_sig000007aa,
      PCIN(18) => blk00000001_sig000007a9,
      PCIN(17) => blk00000001_sig000007a8,
      PCIN(16) => blk00000001_sig000007a7,
      PCIN(15) => blk00000001_sig000007a6,
      PCIN(14) => blk00000001_sig000007a5,
      PCIN(13) => blk00000001_sig000007a4,
      PCIN(12) => blk00000001_sig000007a3,
      PCIN(11) => blk00000001_sig000007a2,
      PCIN(10) => blk00000001_sig000007a1,
      PCIN(9) => blk00000001_sig000007a0,
      PCIN(8) => blk00000001_sig0000079f,
      PCIN(7) => blk00000001_sig0000079e,
      PCIN(6) => blk00000001_sig0000079d,
      PCIN(5) => blk00000001_sig0000079c,
      PCIN(4) => blk00000001_sig0000079b,
      PCIN(3) => blk00000001_sig0000079a,
      PCIN(2) => blk00000001_sig00000799,
      PCIN(1) => blk00000001_sig00000798,
      PCIN(0) => blk00000001_sig00000797,
      ALUMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ALUMODE(1) => blk00000001_sig00000796,
      ALUMODE(0) => blk00000001_sig00000796,
      B(17) => blk00000001_sig000007d7,
      B(16) => blk00000001_sig000007d7,
      B(15) => blk00000001_sig000007d7,
      B(14) => blk00000001_sig000007d6,
      B(13) => blk00000001_sig000007d5,
      B(12) => blk00000001_sig000007d4,
      B(11) => blk00000001_sig000007d3,
      B(10) => blk00000001_sig000007d2,
      B(9) => blk00000001_sig000007d1,
      B(8) => blk00000001_sig000007d0,
      B(7) => blk00000001_sig000007cf,
      B(6) => blk00000001_sig000007ce,
      B(5) => blk00000001_sig000007cd,
      B(4) => blk00000001_sig000007cc,
      B(3) => blk00000001_sig000007cb,
      B(2) => blk00000001_sig000007ca,
      B(1) => blk00000001_sig000007c9,
      B(0) => blk00000001_sig000007c8,
      P(47) => NLW_blk00000001_blk00000d43_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk00000d43_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk00000d43_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk00000d43_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk00000d43_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk00000d43_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk00000d43_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk00000d43_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk00000d43_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk00000d43_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk00000d43_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk00000d43_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk00000d43_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk00000d43_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk00000d43_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk00000d43_P_32_UNCONNECTED,
      P(31) => blk00000001_sig00000755,
      P(30) => blk00000001_sig00000754,
      P(29) => blk00000001_sig00000753,
      P(28) => blk00000001_sig00000752,
      P(27) => blk00000001_sig00000751,
      P(26) => blk00000001_sig00000750,
      P(25) => blk00000001_sig0000074f,
      P(24) => blk00000001_sig0000074e,
      P(23) => blk00000001_sig0000074d,
      P(22) => blk00000001_sig0000074c,
      P(21) => blk00000001_sig0000074b,
      P(20) => blk00000001_sig0000074a,
      P(19) => blk00000001_sig00000749,
      P(18) => blk00000001_sig00000748,
      P(17) => blk00000001_sig00000747,
      P(16) => blk00000001_sig00000746,
      P(15) => blk00000001_sig00000745,
      P(14) => blk00000001_sig00000744,
      P(13) => blk00000001_sig00000743,
      P(12) => blk00000001_sig00000742,
      P(11) => NLW_blk00000001_blk00000d43_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk00000d43_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk00000d43_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk00000d43_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk00000d43_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk00000d43_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk00000d43_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk00000d43_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk00000d43_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk00000d43_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk00000d43_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk00000d43_P_0_UNCONNECTED,
      A(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(24) => blk00000001_sig000007f8,
      A(23) => blk00000001_sig000007f8,
      A(22) => blk00000001_sig000007f8,
      A(21) => blk00000001_sig000007f8,
      A(20) => blk00000001_sig000007f8,
      A(19) => blk00000001_sig000007f8,
      A(18) => blk00000001_sig000007f8,
      A(17) => blk00000001_sig000007f8,
      A(16) => blk00000001_sig000007f8,
      A(15) => blk00000001_sig000007f7,
      A(14) => blk00000001_sig000007f6,
      A(13) => blk00000001_sig000007f5,
      A(12) => blk00000001_sig000007f4,
      A(11) => blk00000001_sig000007f3,
      A(10) => blk00000001_sig000007f2,
      A(9) => blk00000001_sig000007f1,
      A(8) => blk00000001_sig000007f0,
      A(7) => blk00000001_sig000007ef,
      A(6) => blk00000001_sig000007ee,
      A(5) => blk00000001_sig000007ed,
      A(4) => blk00000001_sig000007ec,
      A(3) => blk00000001_sig000007eb,
      A(2) => blk00000001_sig000007ea,
      A(1) => blk00000001_sig000007e9,
      A(0) => blk00000001_sig000007e8,
      PCOUT(47) => NLW_blk00000001_blk00000d43_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk00000d43_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk00000d43_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk00000d43_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk00000d43_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk00000d43_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk00000d43_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk00000d43_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk00000d43_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk00000d43_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk00000d43_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk00000d43_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk00000d43_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk00000d43_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk00000d43_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk00000d43_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk00000d43_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk00000d43_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk00000d43_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk00000d43_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk00000d43_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk00000d43_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk00000d43_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk00000d43_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk00000d43_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk00000d43_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk00000d43_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk00000d43_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk00000d43_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk00000d43_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk00000d43_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk00000d43_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk00000d43_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk00000d43_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk00000d43_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk00000d43_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk00000d43_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk00000d43_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk00000d43_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk00000d43_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk00000d43_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk00000d43_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk00000d43_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk00000d43_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk00000d43_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk00000d43_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk00000d43_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk00000d43_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk00000d43_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk00000d43_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk00000d43_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk00000d43_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk00000d43_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk00000d43_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk00000d43_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk00000d43_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk00000d43_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk00000d43_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk00000d43_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk00000d43_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk00000d43_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk00000d43_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk00000d43_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk00000d43_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk00000d43_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk00000d43_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk00000d43_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk00000d43_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk00000d43_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk00000d43_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk00000d43_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk00000d43_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk00000d43_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk00000d43_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk00000d43_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk00000d43_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk00000d43_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk00000d43_ACOUT_0_UNCONNECTED,
      OPMODE(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(4) => blk00000001_sig000000c0,
      OPMODE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(2) => blk00000001_sig000000c0,
      OPMODE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      OPMODE(0) => blk00000001_sig000000c0,
      CARRYOUT(3) => NLW_blk00000001_blk00000d43_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk00000d43_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk00000d43_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk00000d43_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      BCOUT(17) => NLW_blk00000001_blk00000d43_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk00000d43_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk00000d43_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk00000d43_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk00000d43_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk00000d43_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk00000d43_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk00000d43_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk00000d43_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk00000d43_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk00000d43_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk00000d43_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk00000d43_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk00000d43_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk00000d43_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk00000d43_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk00000d43_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk00000d43_BCOUT_0_UNCONNECTED,
      ACIN(29) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(28) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(27) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(26) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(25) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(24) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(23) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(22) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(21) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(20) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(19) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(18) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(17) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(16) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ACIN(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000fd4,
      Q => blk00000001_sig00000ef5
    );
  blk00000001_blk00000d41 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000efc,
      Q => blk00000001_sig00000fd4,
      Q15 => NLW_blk00000001_blk00000d41_Q15_UNCONNECTED
    );
  blk00000001_blk00000d40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000fd3,
      Q => blk00000001_sig00000ef4
    );
  blk00000001_blk00000d3f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000efd,
      Q => blk00000001_sig00000fd3,
      Q15 => NLW_blk00000001_blk00000d3f_Q15_UNCONNECTED
    );
  blk00000001_blk00000d3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000fd2,
      Q => blk00000001_sig00000ef2
    );
  blk00000001_blk00000d3d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000eff,
      Q => blk00000001_sig00000fd2,
      Q15 => NLW_blk00000001_blk00000d3d_Q15_UNCONNECTED
    );
  blk00000001_blk00000d3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000fd1,
      Q => blk00000001_sig00000e15
    );
  blk00000001_blk00000d3b : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000e22,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_sig00000fd1,
      Q31 => NLW_blk00000001_blk00000d3b_Q31_UNCONNECTED,
      A(4) => blk00000001_sig000000c0,
      A(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A(1) => blk00000001_sig000000c0,
      A(0) => blk00000001_sig000000c0
    );
  blk00000001_blk00000d3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000fd0,
      Q => blk00000001_sig00000ef3
    );
  blk00000001_blk00000d39 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000efe,
      Q => blk00000001_sig00000fd0,
      Q15 => NLW_blk00000001_blk00000d39_Q15_UNCONNECTED
    );
  blk00000001_blk00000d38 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000008e,
      ENBWREN => blk00000001_sig0000008e,
      REGCEAREGCE => blk00000001_sig0000008e,
      REGCEB => blk00000001_sig0000008e,
      RSTRAMARSTRAM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTRAMB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGARSTREG => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(8) => blk00000001_sig00000dbf,
      ADDRARDADDR(7) => blk00000001_sig00000dbe,
      ADDRARDADDR(6) => blk00000001_sig00000dbd,
      ADDRARDADDR(5) => blk00000001_sig00000dbc,
      ADDRARDADDR(4) => blk00000001_sig00000dbb,
      ADDRARDADDR(3) => blk00000001_sig000000c0,
      ADDRARDADDR(2) => blk00000001_sig000000c0,
      ADDRARDADDR(1) => blk00000001_sig000000c0,
      ADDRARDADDR(0) => blk00000001_sig000000c0,
      ADDRBWRADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(9) => blk00000001_sig000000c0,
      ADDRBWRADDR(8) => blk00000001_sig00000dbf,
      ADDRBWRADDR(7) => blk00000001_sig00000dbe,
      ADDRBWRADDR(6) => blk00000001_sig00000dbd,
      ADDRBWRADDR(5) => blk00000001_sig00000dbc,
      ADDRBWRADDR(4) => blk00000001_sig00000dbb,
      ADDRBWRADDR(3) => blk00000001_sig000000c0,
      ADDRBWRADDR(2) => blk00000001_sig000000c0,
      ADDRBWRADDR(1) => blk00000001_sig000000c0,
      ADDRBWRADDR(0) => blk00000001_sig000000c0,
      DIADI(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIBDI(15) => NLW_blk00000001_blk00000d38_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk00000d38_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk00000d38_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk00000d38_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk00000d38_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk00000d38_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk00000d38_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk00000d38_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk00000d38_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk00000d38_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk00000d38_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk00000d38_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk00000d38_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk00000d38_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk00000d38_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk00000d38_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPADIP(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPBDIP(1) => NLW_blk00000001_blk00000d38_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk00000d38_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_sig00000f68,
      DOADO(14) => blk00000001_sig00000f67,
      DOADO(13) => blk00000001_sig00000f66,
      DOADO(12) => blk00000001_sig00000f65,
      DOADO(11) => blk00000001_sig00000f64,
      DOADO(10) => blk00000001_sig00000f63,
      DOADO(9) => blk00000001_sig00000f62,
      DOADO(8) => blk00000001_sig00000f61,
      DOADO(7) => blk00000001_sig00000f60,
      DOADO(6) => blk00000001_sig00000f5f,
      DOADO(5) => blk00000001_sig00000f5e,
      DOADO(4) => blk00000001_sig00000f5d,
      DOADO(3) => blk00000001_sig00000f5c,
      DOADO(2) => blk00000001_sig00000f5b,
      DOADO(1) => blk00000001_sig00000f5a,
      DOADO(0) => blk00000001_sig00000f59,
      DOBDO(15) => blk00000001_sig00000f57,
      DOBDO(14) => blk00000001_sig00000f56,
      DOBDO(13) => blk00000001_sig00000f55,
      DOBDO(12) => blk00000001_sig00000f54,
      DOBDO(11) => blk00000001_sig00000f53,
      DOBDO(10) => blk00000001_sig00000f52,
      DOBDO(9) => blk00000001_sig00000f51,
      DOBDO(8) => blk00000001_sig00000f50,
      DOBDO(7) => blk00000001_sig00000f4f,
      DOBDO(6) => blk00000001_sig00000f4e,
      DOBDO(5) => blk00000001_sig00000f4d,
      DOBDO(4) => blk00000001_sig00000f4c,
      DOBDO(3) => blk00000001_sig00000f4b,
      DOBDO(2) => blk00000001_sig00000f4a,
      DOBDO(1) => blk00000001_sig00000f49,
      DOBDO(0) => blk00000001_sig00000f48,
      DOPADOP(1) => NLW_blk00000001_blk00000d38_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_sig00000f69,
      DOPBDOP(1) => NLW_blk00000001_blk00000d38_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_sig00000f58,
      WEA(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEA(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d37 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000008e,
      ENBWREN => blk00000001_sig0000008e,
      REGCEAREGCE => blk00000001_sig0000008e,
      REGCEB => blk00000001_sig0000008e,
      RSTRAMARSTRAM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTRAMB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGARSTREG => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(8) => blk00000001_sig00000dc4,
      ADDRARDADDR(7) => blk00000001_sig00000dc3,
      ADDRARDADDR(6) => blk00000001_sig00000dc2,
      ADDRARDADDR(5) => blk00000001_sig00000dc1,
      ADDRARDADDR(4) => blk00000001_sig00000dc0,
      ADDRARDADDR(3) => blk00000001_sig000000c0,
      ADDRARDADDR(2) => blk00000001_sig000000c0,
      ADDRARDADDR(1) => blk00000001_sig000000c0,
      ADDRARDADDR(0) => blk00000001_sig000000c0,
      ADDRBWRADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(9) => blk00000001_sig000000c0,
      ADDRBWRADDR(8) => blk00000001_sig00000dc4,
      ADDRBWRADDR(7) => blk00000001_sig00000dc3,
      ADDRBWRADDR(6) => blk00000001_sig00000dc2,
      ADDRBWRADDR(5) => blk00000001_sig00000dc1,
      ADDRBWRADDR(4) => blk00000001_sig00000dc0,
      ADDRBWRADDR(3) => blk00000001_sig000000c0,
      ADDRBWRADDR(2) => blk00000001_sig000000c0,
      ADDRBWRADDR(1) => blk00000001_sig000000c0,
      ADDRBWRADDR(0) => blk00000001_sig000000c0,
      DIADI(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIBDI(15) => NLW_blk00000001_blk00000d37_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk00000d37_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk00000d37_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk00000d37_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk00000d37_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk00000d37_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk00000d37_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk00000d37_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk00000d37_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk00000d37_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk00000d37_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk00000d37_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk00000d37_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk00000d37_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk00000d37_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk00000d37_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPADIP(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPBDIP(1) => NLW_blk00000001_blk00000d37_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk00000d37_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_sig00000f46,
      DOADO(14) => blk00000001_sig00000f45,
      DOADO(13) => blk00000001_sig00000f44,
      DOADO(12) => blk00000001_sig00000f43,
      DOADO(11) => blk00000001_sig00000f42,
      DOADO(10) => blk00000001_sig00000f41,
      DOADO(9) => blk00000001_sig00000f40,
      DOADO(8) => blk00000001_sig00000f3f,
      DOADO(7) => blk00000001_sig00000f3e,
      DOADO(6) => blk00000001_sig00000f3d,
      DOADO(5) => blk00000001_sig00000f3c,
      DOADO(4) => blk00000001_sig00000f3b,
      DOADO(3) => blk00000001_sig00000f3a,
      DOADO(2) => blk00000001_sig00000f39,
      DOADO(1) => blk00000001_sig00000f38,
      DOADO(0) => blk00000001_sig00000f37,
      DOBDO(15) => blk00000001_sig00000f35,
      DOBDO(14) => blk00000001_sig00000f34,
      DOBDO(13) => blk00000001_sig00000f33,
      DOBDO(12) => blk00000001_sig00000f32,
      DOBDO(11) => blk00000001_sig00000f31,
      DOBDO(10) => blk00000001_sig00000f30,
      DOBDO(9) => blk00000001_sig00000f2f,
      DOBDO(8) => blk00000001_sig00000f2e,
      DOBDO(7) => blk00000001_sig00000f2d,
      DOBDO(6) => blk00000001_sig00000f2c,
      DOBDO(5) => blk00000001_sig00000f2b,
      DOBDO(4) => blk00000001_sig00000f2a,
      DOBDO(3) => blk00000001_sig00000f29,
      DOBDO(2) => blk00000001_sig00000f28,
      DOBDO(1) => blk00000001_sig00000f27,
      DOBDO(0) => blk00000001_sig00000f26,
      DOPADOP(1) => NLW_blk00000001_blk00000d37_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_sig00000f47,
      DOPBDOP(1) => NLW_blk00000001_blk00000d37_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_sig00000f36,
      WEA(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEA(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d36 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000008e,
      ENBWREN => blk00000001_sig0000008e,
      REGCEAREGCE => blk00000001_sig0000008e,
      REGCEB => blk00000001_sig0000008e,
      RSTRAMARSTRAM => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTRAMB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGARSTREG => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      RSTREGB => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRARDADDR(8) => blk00000001_sig00000dc9,
      ADDRARDADDR(7) => blk00000001_sig00000dc8,
      ADDRARDADDR(6) => blk00000001_sig00000dc7,
      ADDRARDADDR(5) => blk00000001_sig00000dc6,
      ADDRARDADDR(4) => blk00000001_sig00000dc5,
      ADDRARDADDR(3) => blk00000001_sig000000c0,
      ADDRARDADDR(2) => blk00000001_sig000000c0,
      ADDRARDADDR(1) => blk00000001_sig000000c0,
      ADDRARDADDR(0) => blk00000001_sig000000c0,
      ADDRBWRADDR(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      ADDRBWRADDR(9) => blk00000001_sig000000c0,
      ADDRBWRADDR(8) => blk00000001_sig00000dc9,
      ADDRBWRADDR(7) => blk00000001_sig00000dc8,
      ADDRBWRADDR(6) => blk00000001_sig00000dc7,
      ADDRBWRADDR(5) => blk00000001_sig00000dc6,
      ADDRBWRADDR(4) => blk00000001_sig00000dc5,
      ADDRBWRADDR(3) => blk00000001_sig000000c0,
      ADDRBWRADDR(2) => blk00000001_sig000000c0,
      ADDRBWRADDR(1) => blk00000001_sig000000c0,
      ADDRBWRADDR(0) => blk00000001_sig000000c0,
      DIADI(15) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(14) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(13) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(12) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(11) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(10) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(9) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(8) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(7) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(6) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(5) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(4) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIADI(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIBDI(15) => NLW_blk00000001_blk00000d36_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk00000d36_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk00000d36_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk00000d36_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk00000d36_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk00000d36_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk00000d36_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk00000d36_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk00000d36_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk00000d36_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk00000d36_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk00000d36_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk00000d36_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk00000d36_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk00000d36_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk00000d36_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPADIP(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      DIPBDIP(1) => NLW_blk00000001_blk00000d36_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk00000d36_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_sig00000f24,
      DOADO(14) => blk00000001_sig00000f23,
      DOADO(13) => blk00000001_sig00000f22,
      DOADO(12) => blk00000001_sig00000f21,
      DOADO(11) => blk00000001_sig00000f20,
      DOADO(10) => blk00000001_sig00000f1f,
      DOADO(9) => blk00000001_sig00000f1e,
      DOADO(8) => blk00000001_sig00000f1d,
      DOADO(7) => blk00000001_sig00000f1c,
      DOADO(6) => blk00000001_sig00000f1b,
      DOADO(5) => blk00000001_sig00000f1a,
      DOADO(4) => blk00000001_sig00000f19,
      DOADO(3) => blk00000001_sig00000f18,
      DOADO(2) => blk00000001_sig00000f17,
      DOADO(1) => blk00000001_sig00000f16,
      DOADO(0) => blk00000001_sig00000f15,
      DOBDO(15) => blk00000001_sig00000f13,
      DOBDO(14) => blk00000001_sig00000f12,
      DOBDO(13) => blk00000001_sig00000f11,
      DOBDO(12) => blk00000001_sig00000f10,
      DOBDO(11) => blk00000001_sig00000f0f,
      DOBDO(10) => blk00000001_sig00000f0e,
      DOBDO(9) => blk00000001_sig00000f0d,
      DOBDO(8) => blk00000001_sig00000f0c,
      DOBDO(7) => blk00000001_sig00000f0b,
      DOBDO(6) => blk00000001_sig00000f0a,
      DOBDO(5) => blk00000001_sig00000f09,
      DOBDO(4) => blk00000001_sig00000f08,
      DOBDO(3) => blk00000001_sig00000f07,
      DOBDO(2) => blk00000001_sig00000f06,
      DOBDO(1) => blk00000001_sig00000f05,
      DOBDO(0) => blk00000001_sig00000f04,
      DOPADOP(1) => NLW_blk00000001_blk00000d36_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_sig00000f25,
      DOPBDOP(1) => NLW_blk00000001_blk00000d36_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_sig00000f14,
      WEA(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEA(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(3) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(2) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(1) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      WEBWE(0) => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000d35 : LUT6
    generic map(
      INIT => X"FFFFFFFF22202020"
    )
    port map (
      I0 => blk00000001_sig000000e1,
      I1 => blk00000001_sig000000c3,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig000000c5,
      I4 => blk00000001_sig000000df,
      I5 => blk00000001_sig00000f9e,
      O => blk00000001_sig00000fcf
    );
  blk00000001_blk00000d34 : LUT5
    generic map(
      INIT => X"88888000"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig00000fa0,
      I2 => blk00000001_sig000000df,
      I3 => blk00000001_sig000000c5,
      I4 => blk00000001_sig000000bb,
      O => blk00000001_sig00000fce
    );
  blk00000001_blk00000d33 : MUXF7
    port map (
      I0 => blk00000001_sig00000fce,
      I1 => blk00000001_sig00000fcf,
      S => blk00000001_sig000000ed,
      O => blk00000001_sig00000f83
    );
  blk00000001_blk00000d32 : LUT6
    generic map(
      INIT => X"1515151510101000"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000e1f,
      I4 => blk00000001_sig00000e13,
      I5 => blk00000001_sig000000bb,
      O => blk00000001_sig00000fcd
    );
  blk00000001_blk00000d31 : LUT4
    generic map(
      INIT => X"0444"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig00000e26,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000fcc
    );
  blk00000001_blk00000d30 : MUXF7
    port map (
      I0 => blk00000001_sig00000fcc,
      I1 => blk00000001_sig00000fcd,
      S => blk00000001_sig0000008a,
      O => blk00000001_sig00000f93
    );
  blk00000001_blk00000d2f : INV
    port map (
      I => blk00000001_sig00000b9e,
      O => blk00000001_sig00000b9f
    );
  blk00000001_blk00000d2e : INV
    port map (
      I => blk00000001_sig00000ba0,
      O => blk00000001_sig00000c01
    );
  blk00000001_blk00000d2d : INV
    port map (
      I => blk00000001_sig000008ae,
      O => blk00000001_sig0000087d
    );
  blk00000001_blk00000d2c : INV
    port map (
      I => blk00000001_sig000007c7,
      O => blk00000001_sig0000080a
    );
  blk00000001_blk00000d2b : INV
    port map (
      I => blk00000001_sig000007c7,
      O => blk00000001_sig00000796
    );
  blk00000001_blk00000d2a : INV
    port map (
      I => aresetn,
      O => blk00000001_sig000000cc
    );
  blk00000001_blk00000d29 : FDR
    port map (
      C => aclk,
      D => blk00000001_sig000000cf,
      R => blk00000001_sig000000cc,
      Q => blk00000001_sig00000fcb
    );
  blk00000001_blk00000d28 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000015b,
      I2 => blk00000001_sig0000017e,
      O => blk00000001_sig00000fca
    );
  blk00000001_blk00000d27 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000015a,
      I2 => blk00000001_sig0000017d,
      O => blk00000001_sig00000fc9
    );
  blk00000001_blk00000d26 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000159,
      I2 => blk00000001_sig0000017c,
      O => blk00000001_sig00000fc8
    );
  blk00000001_blk00000d25 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000158,
      I2 => blk00000001_sig0000017b,
      O => blk00000001_sig00000fc7
    );
  blk00000001_blk00000d24 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000157,
      I2 => blk00000001_sig0000017a,
      O => blk00000001_sig00000fc6
    );
  blk00000001_blk00000d23 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000156,
      I2 => blk00000001_sig00000179,
      O => blk00000001_sig00000fc5
    );
  blk00000001_blk00000d22 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000155,
      I2 => blk00000001_sig00000178,
      O => blk00000001_sig00000fc4
    );
  blk00000001_blk00000d21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000154,
      I2 => blk00000001_sig00000177,
      O => blk00000001_sig00000fc3
    );
  blk00000001_blk00000d20 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000153,
      I2 => blk00000001_sig00000176,
      O => blk00000001_sig00000fc2
    );
  blk00000001_blk00000d1f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000152,
      I2 => blk00000001_sig00000175,
      O => blk00000001_sig00000fc1
    );
  blk00000001_blk00000d1e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000151,
      I2 => blk00000001_sig00000174,
      O => blk00000001_sig00000fc0
    );
  blk00000001_blk00000d1d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000150,
      I2 => blk00000001_sig00000173,
      O => blk00000001_sig00000fbf
    );
  blk00000001_blk00000d1c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014f,
      I2 => blk00000001_sig00000172,
      O => blk00000001_sig00000fbe
    );
  blk00000001_blk00000d1b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014e,
      I2 => blk00000001_sig00000171,
      O => blk00000001_sig00000fbd
    );
  blk00000001_blk00000d1a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014d,
      I2 => blk00000001_sig00000170,
      O => blk00000001_sig00000fbc
    );
  blk00000001_blk00000d19 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014c,
      I2 => blk00000001_sig0000016f,
      O => blk00000001_sig00000fbb
    );
  blk00000001_blk00000d18 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014b,
      I2 => blk00000001_sig0000016e,
      O => blk00000001_sig00000fba
    );
  blk00000001_blk00000d17 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000014a,
      I2 => blk00000001_sig0000016d,
      O => blk00000001_sig00000fb9
    );
  blk00000001_blk00000d16 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000149,
      I2 => blk00000001_sig0000016c,
      O => blk00000001_sig00000fb8
    );
  blk00000001_blk00000d15 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000148,
      I2 => blk00000001_sig0000016b,
      O => blk00000001_sig00000fb7
    );
  blk00000001_blk00000d14 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000147,
      I2 => blk00000001_sig0000016a,
      O => blk00000001_sig00000fb6
    );
  blk00000001_blk00000d13 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000146,
      I2 => blk00000001_sig00000169,
      O => blk00000001_sig00000fb5
    );
  blk00000001_blk00000d12 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000145,
      I2 => blk00000001_sig00000168,
      O => blk00000001_sig00000fb4
    );
  blk00000001_blk00000d11 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000144,
      I2 => blk00000001_sig00000167,
      O => blk00000001_sig00000fb3
    );
  blk00000001_blk00000d10 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000143,
      I2 => blk00000001_sig00000166,
      O => blk00000001_sig00000fb2
    );
  blk00000001_blk00000d0f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000142,
      I2 => blk00000001_sig00000165,
      O => blk00000001_sig00000fb1
    );
  blk00000001_blk00000d0e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000141,
      I2 => blk00000001_sig00000164,
      O => blk00000001_sig00000fb0
    );
  blk00000001_blk00000d0d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig00000140,
      I2 => blk00000001_sig00000163,
      O => blk00000001_sig00000faf
    );
  blk00000001_blk00000d0c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000013f,
      I2 => blk00000001_sig00000162,
      O => blk00000001_sig00000fae
    );
  blk00000001_blk00000d0b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000013e,
      I2 => blk00000001_sig00000161,
      O => blk00000001_sig00000fad
    );
  blk00000001_blk00000d0a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000013d,
      I2 => blk00000001_sig00000160,
      O => blk00000001_sig00000fac
    );
  blk00000001_blk00000d09 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000013c,
      I2 => blk00000001_sig0000015f,
      O => blk00000001_sig00000fab
    );
  blk00000001_blk00000d08 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000fa8,
      I1 => blk00000001_sig0000013b,
      I2 => blk00000001_sig0000015e,
      O => blk00000001_sig00000faa
    );
  blk00000001_blk00000d07 : LUT4
    generic map(
      INIT => X"FBFF"
    )
    port map (
      I0 => blk00000001_sig000000f3,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig000000f8,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000fa9
    );
  blk00000001_blk00000d06 : LUT3
    generic map(
      INIT => X"20"
    )
    port map (
      I0 => blk00000001_sig0000015c,
      I1 => blk00000001_sig0000013a,
      I2 => blk00000001_sig00000101,
      O => blk00000001_sig00000fa8
    );
  blk00000001_blk00000d05 : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000de8,
      I2 => blk00000001_sig00000e22,
      O => blk00000001_sig00000da5
    );
  blk00000001_blk00000d04 : LUT4
    generic map(
      INIT => X"1F0C"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig0000008d,
      I2 => blk00000001_sig00000e15,
      I3 => blk00000001_sig00000e22,
      O => blk00000001_sig00000f91
    );
  blk00000001_blk00000d03 : LUT4
    generic map(
      INIT => X"1F0C"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig0000008d,
      I2 => blk00000001_sig00000e20,
      I3 => blk00000001_sig00000e21,
      O => blk00000001_sig00000f90
    );
  blk00000001_blk00000d02 : LUT6
    generic map(
      INIT => X"FFFFFFFF80888080"
    )
    port map (
      I0 => blk00000001_sig00000dea,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig000001a8,
      I3 => blk00000001_sig0000008d,
      I4 => blk00000001_sig00000e12,
      I5 => blk00000001_sig000001b2,
      O => blk00000001_sig00000e6c
    );
  blk00000001_blk00000d01 : LUT5
    generic map(
      INIT => X"AAEAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000e62,
      I1 => blk00000001_sig000000bc,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000e1e,
      I4 => blk00000001_sig000001a8,
      O => blk00000001_sig00000e5d
    );
  blk00000001_blk00000d00 : LUT5
    generic map(
      INIT => X"EAAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000df2,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig00000e25,
      O => blk00000001_sig00000e4e
    );
  blk00000001_blk00000cff : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig0000008f,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000e26,
      O => blk00000001_sig00000e41
    );
  blk00000001_blk00000cfe : LUT6
    generic map(
      INIT => X"40404040404040EF"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_event_tlast_missing,
      I2 => blk00000001_sig000000ec,
      I3 => blk00000001_sig00000102,
      I4 => blk00000001_sig000000c3,
      I5 => blk00000001_sig000000c5,
      O => blk00000001_sig00000f88
    );
  blk00000001_blk00000cfd : LUT6
    generic map(
      INIT => X"EE6ECC6CEEEEECEC"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig000000f8,
      I4 => blk00000001_sig000000c4,
      I5 => blk00000001_sig000000f4,
      O => blk00000001_sig00000f80
    );
  blk00000001_blk00000cfc : LUT6
    generic map(
      INIT => X"44444444444F4444"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000ec,
      I2 => blk00000001_sig00000102,
      I3 => blk00000001_sig000000f3,
      I4 => blk00000001_sig0000008e,
      I5 => blk00000001_sig000000c5,
      O => blk00000001_sig00000f82
    );
  blk00000001_blk00000cfb : LUT3
    generic map(
      INIT => X"02"
    )
    port map (
      I0 => blk00000001_sig0000008b,
      I1 => blk00000001_sig000000e3,
      I2 => blk00000001_sig000000f8,
      O => blk00000001_sig00000f8b
    );
  blk00000001_blk00000cfa : LUT5
    generic map(
      INIT => X"555D0008"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig000000f3,
      I3 => blk00000001_sig00000101,
      I4 => NlwRenamedSig_OI_event_data_in_channel_halt,
      O => blk00000001_sig00000f87
    );
  blk00000001_blk00000cf9 : LUT6
    generic map(
      INIT => X"5410101010101010"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig00000e13,
      I3 => blk00000001_sig00000e24,
      I4 => blk00000001_sig000000bc,
      I5 => blk00000001_sig00000dea,
      O => blk00000001_sig00000f9c
    );
  blk00000001_blk00000cf8 : LUT6
    generic map(
      INIT => X"0111010100100000"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e22,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig000001a7,
      I4 => blk00000001_sig000002e2,
      I5 => blk00000001_sig000000bf,
      O => blk00000001_sig00000f98
    );
  blk00000001_blk00000cf7 : LUT4
    generic map(
      INIT => X"5540"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig000000bc,
      I3 => blk00000001_sig00000e16,
      O => blk00000001_sig00000f8d
    );
  blk00000001_blk00000cf6 : LUT5
    generic map(
      INIT => X"15151000"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e0f,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000e12,
      I4 => blk00000001_sig000000bc,
      O => blk00000001_sig00000f92
    );
  blk00000001_blk00000cf5 : LUT4
    generic map(
      INIT => X"BA10"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => blk00000001_sig0000008b,
      I2 => blk00000001_sig000000fd,
      I3 => blk00000001_sig000000f7,
      O => blk00000001_sig00000f8a
    );
  blk00000001_blk00000cf4 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig00000e27,
      I4 => blk00000001_sig00000e12,
      O => blk00000001_sig00000f9b
    );
  blk00000001_blk00000cf3 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig00000e24,
      I3 => blk00000001_sig00000dea,
      I4 => blk00000001_sig000000bd,
      O => blk00000001_sig00000f9a
    );
  blk00000001_blk00000cf2 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => aclken,
      I2 => blk00000001_sig000000ff,
      I3 => blk00000001_sig000000be,
      I4 => NlwRenamedSig_OI_event_data_out_channel_halt,
      O => blk00000001_sig00000f97
    );
  blk00000001_blk00000cf1 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => aclken,
      I2 => blk00000001_sig00000100,
      I3 => blk00000001_sig000000fa,
      I4 => NlwRenamedSig_OI_event_status_channel_halt,
      O => blk00000001_sig00000f96
    );
  blk00000001_blk00000cf0 : LUT5
    generic map(
      INIT => X"11510040"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => blk00000001_sig0000008e,
      I2 => blk00000001_sig000000de,
      I3 => blk00000001_sig000000be,
      I4 => blk00000001_sig000000dd,
      O => blk00000001_sig00000f95
    );
  blk00000001_blk00000cef : LUT6
    generic map(
      INIT => X"5410101010101010"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_event_fft_overflow,
      I3 => m_axis_data_tready,
      I4 => NlwRenamedSig_OI_m_axis_data_tuser_8_Q,
      I5 => NlwRenamedSig_OI_m_axis_data_tvalid,
      O => blk00000001_sig00000f94
    );
  blk00000001_blk00000cee : LUT6
    generic map(
      INIT => X"0454044404440444"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig000002e2,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig000001a9,
      I4 => blk00000001_sig000001aa,
      I5 => blk00000001_sig00000367,
      O => blk00000001_sig00000f99
    );
  blk00000001_blk00000ced : LUT5
    generic map(
      INIT => X"FFFF5C4C"
    )
    port map (
      I0 => blk00000001_sig00000e25,
      I1 => blk00000001_sig00000e1e,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig000001a8,
      I4 => blk00000001_sig0000008d,
      O => blk00000001_sig00000f8e
    );
  blk00000001_blk00000cec : LUT6
    generic map(
      INIT => X"FFFFFFFFBAAA8AAA"
    )
    port map (
      I0 => blk00000001_sig000000f1,
      I1 => blk00000001_sig000000f8,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig000000ca,
      I5 => blk00000001_sig000000d7,
      O => blk00000001_sig00000f7a
    );
  blk00000001_blk00000ceb : LUT6
    generic map(
      INIT => X"AAAAAACAAAAAAAAA"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => blk00000001_sig000000bf,
      I2 => blk00000001_sig000000c6,
      I3 => blk00000001_sig000000f8,
      I4 => blk00000001_sig00000fa7,
      I5 => blk00000001_sig000000c4,
      O => blk00000001_sig00000f8c
    );
  blk00000001_blk00000cea : LUT2
    generic map(
      INIT => X"D"
    )
    port map (
      I0 => blk00000001_sig000000be,
      I1 => blk00000001_sig000000eb,
      O => blk00000001_sig00000fa7
    );
  blk00000001_blk00000ce9 : LUT6
    generic map(
      INIT => X"FFFFFFFFAAA9AAAA"
    )
    port map (
      I0 => blk00000001_sig000000f0,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000ee,
      I3 => blk00000001_sig000000ef,
      I4 => blk00000001_sig000000da,
      I5 => blk00000001_sig000000d7,
      O => blk00000001_sig00000f7b
    );
  blk00000001_blk00000ce8 : LUT6
    generic map(
      INIT => X"FFFFFFFFBAAA8AAA"
    )
    port map (
      I0 => blk00000001_sig000000f2,
      I1 => blk00000001_sig000000f8,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig000000c9,
      I5 => blk00000001_sig000000d7,
      O => blk00000001_sig00000f79
    );
  blk00000001_blk00000ce7 : LUT6
    generic map(
      INIT => X"FFFF7300FFFF5000"
    )
    port map (
      I0 => blk00000001_sig000000f4,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig00000f7e,
      I5 => blk00000001_sig000000c4,
      O => blk00000001_sig00000f7f
    );
  blk00000001_blk00000ce6 : LUT6
    generic map(
      INIT => X"FFFF7300FFFF5000"
    )
    port map (
      I0 => blk00000001_sig000000f4,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig00000f7c,
      I5 => blk00000001_sig000000c4,
      O => blk00000001_sig00000f7d
    );
  blk00000001_blk00000ce5 : LUT6
    generic map(
      INIT => X"ECECEEECCCCCCCCC"
    )
    port map (
      I0 => blk00000001_sig00000dea,
      I1 => blk00000001_sig000001b1,
      I2 => blk00000001_sig000001a8,
      I3 => blk00000001_sig00000e12,
      I4 => blk00000001_sig0000008d,
      I5 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e6b
    );
  blk00000001_blk00000ce4 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000e61,
      I1 => blk00000001_sig000001a8,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e5c
    );
  blk00000001_blk00000ce3 : LUT5
    generic map(
      INIT => X"ECCCCCCC"
    )
    port map (
      I0 => blk00000001_sig00000e25,
      I1 => blk00000001_sig00000df1,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e4d
    );
  blk00000001_blk00000ce2 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig00000090,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e40
    );
  blk00000001_blk00000ce1 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000e60,
      I1 => blk00000001_sig000001a8,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e5b
    );
  blk00000001_blk00000ce0 : LUT5
    generic map(
      INIT => X"ECCCCCCC"
    )
    port map (
      I0 => blk00000001_sig00000e25,
      I1 => blk00000001_sig00000df0,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e4c
    );
  blk00000001_blk00000cdf : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig00000091,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e3f
    );
  blk00000001_blk00000cde : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000e5f,
      I1 => blk00000001_sig000001a8,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e5a
    );
  blk00000001_blk00000cdd : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig00000092,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e3e
    );
  blk00000001_blk00000cdc : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig00000093,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e3d
    );
  blk00000001_blk00000cdb : LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      I0 => blk00000001_sig000000e1,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig000000df,
      I3 => blk00000001_sig000000c5,
      O => blk00000001_sig000000d5
    );
  blk00000001_blk00000cda : LUT5
    generic map(
      INIT => X"0040AAEA"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000101,
      I2 => blk00000001_sig0000015c,
      I3 => blk00000001_sig000000dc,
      I4 => blk00000001_sig00000117,
      O => blk00000001_sig00000f86
    );
  blk00000001_blk00000cd9 : LUT6
    generic map(
      INIT => X"FFFF0CCCFFFF0C4C"
    )
    port map (
      I0 => blk00000001_sig000000df,
      I1 => blk00000001_sig000000f3,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000fa6,
      I4 => blk00000001_sig000000d6,
      I5 => blk00000001_sig000000c5,
      O => blk00000001_sig00000f84
    );
  blk00000001_blk00000cd8 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig000000be,
      I1 => blk00000001_sig000000de,
      O => blk00000001_sig00000fa6
    );
  blk00000001_blk00000cd7 : LUT6
    generic map(
      INIT => X"FFFFFFFFAAAAAA2A"
    )
    port map (
      I0 => blk00000001_sig00000101,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig000000f8,
      I4 => blk00000001_sig000000f3,
      I5 => blk00000001_sig00000116,
      O => blk00000001_sig00000f85
    );
  blk00000001_blk00000cd6 : LUT6
    generic map(
      INIT => X"FFFFFFFFFFFFFFFE"
    )
    port map (
      I0 => blk00000001_sig00000f72,
      I1 => blk00000001_sig00000f74,
      I2 => blk00000001_sig00000fa5,
      I3 => blk00000001_sig00000f9f,
      I4 => blk00000001_sig00000f71,
      I5 => blk00000001_sig00000f78,
      O => blk00000001_sig00000c8a
    );
  blk00000001_blk00000cd5 : LUT5
    generic map(
      INIT => X"FFFF7FFE"
    )
    port map (
      I0 => blk00000001_sig00000397,
      I1 => blk00000001_sig000006ce,
      I2 => blk00000001_sig000006cd,
      I3 => blk00000001_sig000006cc,
      I4 => blk00000001_sig00000f73,
      O => blk00000001_sig00000fa5
    );
  blk00000001_blk00000cd4 : LUT5
    generic map(
      INIT => X"AA9AAAAA"
    )
    port map (
      I0 => blk00000001_sig000000ee,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig000000f8,
      I4 => blk00000001_sig0000008e,
      O => blk00000001_sig00000f7e
    );
  blk00000001_blk00000cd3 : LUT6
    generic map(
      INIT => X"AAAAA9AAAAAAAAAA"
    )
    port map (
      I0 => blk00000001_sig000000ef,
      I1 => blk00000001_sig000000ee,
      I2 => blk00000001_sig000000c6,
      I3 => blk00000001_sig000000be,
      I4 => blk00000001_sig000000f8,
      I5 => blk00000001_sig0000008e,
      O => blk00000001_sig00000f7c
    );
  blk00000001_blk00000cd2 : LUT5
    generic map(
      INIT => X"40EA00AA"
    )
    port map (
      I0 => blk00000001_sig000000eb,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig000000cb,
      I4 => blk00000001_sig000000c4,
      O => blk00000001_sig00000f81
    );
  blk00000001_blk00000cd1 : LUT5
    generic map(
      INIT => X"F0FCFEFC"
    )
    port map (
      I0 => blk00000001_sig00000e14,
      I1 => blk00000001_sig00000e1f,
      I2 => blk00000001_sig0000008d,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig0000008a,
      O => blk00000001_sig00000f8f
    );
  blk00000001_blk00000cd0 : LUT6
    generic map(
      INIT => X"FFF4FFFEFFF5FFFF"
    )
    port map (
      I0 => blk00000001_sig000006dd,
      I1 => blk00000001_sig000003e7,
      I2 => blk00000001_sig00000f77,
      I3 => blk00000001_sig00000f76,
      I4 => blk00000001_sig00000fa4,
      I5 => blk00000001_sig00000fa3,
      O => blk00000001_sig00000f78
    );
  blk00000001_blk00000ccf : LUT4
    generic map(
      INIT => X"AAAB"
    )
    port map (
      I0 => blk00000001_sig000006d7,
      I1 => blk00000001_sig000006d5,
      I2 => blk00000001_sig000006d6,
      I3 => blk00000001_sig000003c7,
      O => blk00000001_sig00000fa4
    );
  blk00000001_blk00000cce : LUT6
    generic map(
      INIT => X"1010101010101011"
    )
    port map (
      I0 => blk00000001_sig000006dc,
      I1 => blk00000001_sig000006db,
      I2 => blk00000001_sig000006d7,
      I3 => blk00000001_sig000003c7,
      I4 => blk00000001_sig000006d6,
      I5 => blk00000001_sig000006d5,
      O => blk00000001_sig00000fa3
    );
  blk00000001_blk00000ccd : LUT6
    generic map(
      INIT => X"FFF7FFF2FFFFFFFA"
    )
    port map (
      I0 => blk00000001_sig000006d4,
      I1 => blk00000001_sig000003b7,
      I2 => blk00000001_sig00000f6f,
      I3 => blk00000001_sig00000f70,
      I4 => blk00000001_sig00000fa1,
      I5 => blk00000001_sig00000fa2,
      O => blk00000001_sig00000f71
    );
  blk00000001_blk00000ccc : LUT6
    generic map(
      INIT => X"8000000088888888"
    )
    port map (
      I0 => blk00000001_sig000006d3,
      I1 => blk00000001_sig000006d2,
      I2 => blk00000001_sig000006d8,
      I3 => blk00000001_sig000003d7,
      I4 => blk00000001_sig000006d9,
      I5 => blk00000001_sig000006da,
      O => blk00000001_sig00000fa2
    );
  blk00000001_blk00000ccb : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_sig000006da,
      I1 => blk00000001_sig000003d7,
      I2 => blk00000001_sig000006d9,
      I3 => blk00000001_sig000006d8,
      O => blk00000001_sig00000fa1
    );
  blk00000001_blk00000cca : LUT4
    generic map(
      INIT => X"F7FF"
    )
    port map (
      I0 => blk00000001_sig00000102,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig000000f3,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000f9d
    );
  blk00000001_blk00000cc9 : LUT6
    generic map(
      INIT => X"00002000AAAAAAAA"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig000000f3,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig000000f8,
      I5 => blk00000001_sig00000101,
      O => blk00000001_sig00000117
    );
  blk00000001_blk00000cc8 : LUT6
    generic map(
      INIT => X"ECECEEECCCCCCCCC"
    )
    port map (
      I0 => blk00000001_sig00000dea,
      I1 => blk00000001_sig000001b0,
      I2 => blk00000001_sig000001a8,
      I3 => blk00000001_sig00000e12,
      I4 => blk00000001_sig0000008d,
      I5 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e6a
    );
  blk00000001_blk00000cc7 : LUT5
    generic map(
      INIT => X"ECCCCCCC"
    )
    port map (
      I0 => blk00000001_sig00000e25,
      I1 => blk00000001_sig00000def,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e4b
    );
  blk00000001_blk00000cc6 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000e5e,
      I1 => blk00000001_sig000001a8,
      I2 => blk00000001_sig00000e1e,
      I3 => blk00000001_sig000000bc,
      I4 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e59
    );
  blk00000001_blk00000cc5 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig00000094,
      I1 => blk00000001_sig00000e26,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000e3c
    );
  blk00000001_blk00000cc4 : LUT6
    generic map(
      INIT => X"0808080008000800"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig000000e1,
      I2 => blk00000001_sig000000f3,
      I3 => blk00000001_sig000000bb,
      I4 => blk00000001_sig000000df,
      I5 => blk00000001_sig000000c5,
      O => blk00000001_sig000000d9
    );
  blk00000001_blk00000cc3 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig000000e1,
      I1 => blk00000001_sig000000f3,
      O => blk00000001_sig00000fa0
    );
  blk00000001_blk00000cc2 : LUT6
    generic map(
      INIT => X"555555554A4AAA4A"
    )
    port map (
      I0 => blk00000001_sig000000fb,
      I1 => blk00000001_sig000000fc,
      I2 => aclken,
      I3 => blk00000001_sig000000c5,
      I4 => blk00000001_sig00000f9d,
      I5 => blk00000001_sig000000c2,
      O => blk00000001_sig000000c8
    );
  blk00000001_blk00000cc1 : LUT6
    generic map(
      INIT => X"77777777AEAEEEAE"
    )
    port map (
      I0 => blk00000001_sig000000fc,
      I1 => blk00000001_sig000000fb,
      I2 => aclken,
      I3 => blk00000001_sig000000c5,
      I4 => blk00000001_sig00000f9d,
      I5 => blk00000001_sig000000c2,
      O => blk00000001_sig000000cd
    );
  blk00000001_blk00000cc0 : LUT6
    generic map(
      INIT => X"3C3C3C3CD0F0D0D0"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000fb,
      I2 => blk00000001_sig000000fc,
      I3 => blk00000001_sig00000f9d,
      I4 => blk00000001_sig000000c5,
      I5 => blk00000001_sig000000c2,
      O => blk00000001_sig000000c7
    );
  blk00000001_blk00000cbf : LUT4
    generic map(
      INIT => X"EF40"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_event_frame_started,
      I2 => blk00000001_sig000000ed,
      I3 => blk00000001_sig000000d9,
      O => blk00000001_sig00000f89
    );
  blk00000001_blk00000cbe : LUT5
    generic map(
      INIT => X"FFFF7FFE"
    )
    port map (
      I0 => blk00000001_sig00000377,
      I1 => blk00000001_sig000006c8,
      I2 => blk00000001_sig000006c7,
      I3 => blk00000001_sig000006c6,
      I4 => blk00000001_sig00000f75,
      O => blk00000001_sig00000f9f
    );
  blk00000001_blk00000cbd : LUT6
    generic map(
      INIT => X"AAAAAAAAAAAAAAA9"
    )
    port map (
      I0 => blk00000001_sig000000f2,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000f0,
      I3 => blk00000001_sig000000ef,
      I4 => blk00000001_sig000000ee,
      I5 => blk00000001_sig000000c6,
      O => blk00000001_sig000000c9
    );
  blk00000001_blk00000cbc : LUT2
    generic map(
      INIT => X"7"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000ed,
      O => blk00000001_sig00000f9e
    );
  blk00000001_blk00000cbb : LUT5
    generic map(
      INIT => X"55755555"
    )
    port map (
      I0 => blk00000001_sig00000101,
      I1 => blk00000001_sig000000f3,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig000000f8,
      I4 => blk00000001_sig00000fcb,
      O => blk00000001_sig00000139
    );
  blk00000001_blk00000cba : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f9c,
      Q => blk00000001_sig00000e13
    );
  blk00000001_blk00000cb9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f9b,
      Q => blk00000001_sig00000e12
    );
  blk00000001_blk00000cb8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f9a,
      Q => blk00000001_sig000000bd
    );
  blk00000001_blk00000cb7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f99,
      Q => blk00000001_sig000002e2
    );
  blk00000001_blk00000cb6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f98,
      Q => blk00000001_sig000000bf
    );
  blk00000001_blk00000cb5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f97,
      Q => NlwRenamedSig_OI_event_data_out_channel_halt
    );
  blk00000001_blk00000cb4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f96,
      Q => NlwRenamedSig_OI_event_status_channel_halt
    );
  blk00000001_blk00000cb3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f95,
      Q => blk00000001_sig000000dd
    );
  blk00000001_blk00000cb2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f94,
      Q => NlwRenamedSig_OI_event_fft_overflow
    );
  blk00000001_blk00000cb1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f93,
      Q => blk00000001_sig000000bb
    );
  blk00000001_blk00000cb0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f92,
      Q => blk00000001_sig000000bc
    );
  blk00000001_blk00000caf : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f91,
      Q => blk00000001_sig00000e22
    );
  blk00000001_blk00000cae : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f90,
      Q => blk00000001_sig00000e21
    );
  blk00000001_blk00000cad : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f8f,
      Q => blk00000001_sig00000e1f
    );
  blk00000001_blk00000cac : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f8e,
      Q => blk00000001_sig00000e1e
    );
  blk00000001_blk00000cab : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f8d,
      Q => blk00000001_sig00000e16
    );
  blk00000001_blk00000caa : FD
    port map (
      C => aclk,
      D => blk00000001_sig00000f8c,
      Q => blk00000001_sig000000f6
    );
  blk00000001_blk00000ca9 : FD
    port map (
      C => aclk,
      D => blk00000001_sig00000f8b,
      Q => blk00000001_sig000000fd
    );
  blk00000001_blk00000ca8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f8a,
      Q => blk00000001_sig000000f7
    );
  blk00000001_blk00000ca7 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f89,
      R => blk00000001_sig000000f8,
      Q => NlwRenamedSig_OI_event_frame_started
    );
  blk00000001_blk00000ca6 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f88,
      R => blk00000001_sig000000f8,
      Q => NlwRenamedSig_OI_event_tlast_missing
    );
  blk00000001_blk00000ca5 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f87,
      R => blk00000001_sig000000f8,
      Q => NlwRenamedSig_OI_event_data_in_channel_halt
    );
  blk00000001_blk00000ca4 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f86,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013a
    );
  blk00000001_blk00000ca3 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f85,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000101
    );
  blk00000001_blk00000ca2 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f84,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f3
    );
  blk00000001_blk00000ca1 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f83,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000ed
    );
  blk00000001_blk00000ca0 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f82,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000ec
    );
  blk00000001_blk00000c9f : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f81,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000eb
    );
  blk00000001_blk00000c9e : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f80,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000c6
    );
  blk00000001_blk00000c9d : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f7f,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000ee
    );
  blk00000001_blk00000c9c : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f7d,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000ef
    );
  blk00000001_blk00000c9b : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f7b,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f0
    );
  blk00000001_blk00000c9a : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f7a,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f1
    );
  blk00000001_blk00000c99 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000f79,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f2
    );
  blk00000001_blk00000c98 : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_sig000006cb,
      I1 => blk00000001_sig000006c9,
      I2 => blk00000001_sig000006ca,
      I3 => blk00000001_sig00000387,
      O => blk00000001_sig00000f77
    );
  blk00000001_blk00000c97 : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_sig000006d4,
      I1 => blk00000001_sig000006d2,
      I2 => blk00000001_sig000006d3,
      I3 => blk00000001_sig000003b7,
      O => blk00000001_sig00000f76
    );
  blk00000001_blk00000c96 : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_sig000006da,
      I1 => blk00000001_sig000006d8,
      I2 => blk00000001_sig000006d9,
      I3 => blk00000001_sig000003d7,
      O => blk00000001_sig00000f75
    );
  blk00000001_blk00000c95 : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_sig000006d1,
      I1 => blk00000001_sig000006cf,
      I2 => blk00000001_sig000006d0,
      I3 => blk00000001_sig000003a7,
      O => blk00000001_sig00000f74
    );
  blk00000001_blk00000c94 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_sig000006cb,
      I1 => blk00000001_sig000006c9,
      I2 => blk00000001_sig000006ca,
      I3 => blk00000001_sig00000387,
      O => blk00000001_sig00000f73
    );
  blk00000001_blk00000c93 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_sig000006d1,
      I1 => blk00000001_sig000006cf,
      I2 => blk00000001_sig000006d0,
      I3 => blk00000001_sig000003a7,
      O => blk00000001_sig00000f72
    );
  blk00000001_blk00000c92 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_sig000006d7,
      I1 => blk00000001_sig000006d5,
      I2 => blk00000001_sig000006d6,
      I3 => blk00000001_sig000003c7,
      O => blk00000001_sig00000f70
    );
  blk00000001_blk00000c91 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_sig000006dd,
      I1 => blk00000001_sig000006db,
      I2 => blk00000001_sig000006dc,
      I3 => blk00000001_sig000003e7,
      O => blk00000001_sig00000f6f
    );
  blk00000001_blk00000c90 : LUT6
    generic map(
      INIT => X"C8C8C0C800000000"
    )
    port map (
      I0 => blk00000001_sig00000101,
      I1 => blk00000001_sig00000f6d,
      I2 => blk00000001_sig00000f6b,
      I3 => blk00000001_sig000000c5,
      I4 => blk00000001_sig00000f6e,
      I5 => blk00000001_sig00000f6c,
      O => blk00000001_sig000000cf
    );
  blk00000001_blk00000c8f : LUT5
    generic map(
      INIT => X"FF8FFFAF"
    )
    port map (
      I0 => blk00000001_sig0000015d,
      I1 => blk00000001_sig0000015c,
      I2 => blk00000001_sig00000101,
      I3 => blk00000001_sig0000013a,
      I4 => blk00000001_sig000000dc,
      O => blk00000001_sig00000f6e
    );
  blk00000001_blk00000c8e : LUT3
    generic map(
      INIT => X"2A"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig00000100,
      I2 => blk00000001_sig000000fa,
      O => blk00000001_sig00000f6d
    );
  blk00000001_blk00000c8d : LUT6
    generic map(
      INIT => X"13111F1F11111F1F"
    )
    port map (
      I0 => blk00000001_sig000000fe,
      I1 => blk00000001_sig000000ff,
      I2 => blk00000001_sig000000bd,
      I3 => blk00000001_sig000000c6,
      I4 => blk00000001_sig000000be,
      I5 => blk00000001_sig000000c4,
      O => blk00000001_sig00000f6c
    );
  blk00000001_blk00000c8c : LUT2
    generic map(
      INIT => X"D"
    )
    port map (
      I0 => blk00000001_sig000000bb,
      I1 => blk00000001_sig000000f3,
      O => blk00000001_sig00000f6b
    );
  blk00000001_blk00000c8b : LUT6
    generic map(
      INIT => X"0000200000000000"
    )
    port map (
      I0 => blk00000001_sig00000102,
      I1 => blk00000001_sig000000f3,
      I2 => blk00000001_sig000000bb,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig00000f6a,
      I5 => blk00000001_sig000000c5,
      O => blk00000001_sig000000c2
    );
  blk00000001_blk00000c8a : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000fc,
      I2 => blk00000001_sig000000fb,
      O => blk00000001_sig00000f6a
    );
  blk00000001_blk00000c89 : LUT4
    generic map(
      INIT => X"9996"
    )
    port map (
      I0 => blk00000001_sig00000df0,
      I1 => blk00000001_sig00000df2,
      I2 => blk00000001_sig00000def,
      I3 => blk00000001_sig00000df1,
      O => blk00000001_sig00000eb9
    );
  blk00000001_blk00000c88 : LUT4
    generic map(
      INIT => X"9996"
    )
    port map (
      I0 => blk00000001_sig00000ea3,
      I1 => blk00000001_sig00000ea5,
      I2 => blk00000001_sig00000ea2,
      I3 => blk00000001_sig00000ea4,
      O => blk00000001_sig00000eb8
    );
  blk00000001_blk00000c87 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000def,
      I1 => blk00000001_sig00000df1,
      O => blk00000001_sig00000eb7
    );
  blk00000001_blk00000c86 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ea2,
      I1 => blk00000001_sig00000ea4,
      O => blk00000001_sig00000eb6
    );
  blk00000001_blk00000c85 : LUT3
    generic map(
      INIT => X"02"
    )
    port map (
      I0 => blk00000001_sig000001b0,
      I1 => blk00000001_sig000001b2,
      I2 => blk00000001_sig000001b1,
      O => blk00000001_sig00000e94
    );
  blk00000001_blk00000c84 : LUT3
    generic map(
      INIT => X"01"
    )
    port map (
      I0 => blk00000001_sig000001b0,
      I1 => blk00000001_sig000001b2,
      I2 => blk00000001_sig000001b1,
      O => blk00000001_sig00000e93
    );
  blk00000001_blk00000c83 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ea7,
      I1 => blk00000001_sig00000ea6,
      O => blk00000001_sig00000e92
    );
  blk00000001_blk00000c82 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_sig00000e97,
      I1 => blk00000001_sig00000e98,
      I2 => blk00000001_sig00000eac,
      O => blk00000001_sig00000e8f
    );
  blk00000001_blk00000c81 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_sig00000e95,
      I1 => blk00000001_sig00000e96,
      I2 => blk00000001_sig00000eab,
      O => blk00000001_sig00000e8e
    );
  blk00000001_blk00000c80 : LUT4
    generic map(
      INIT => X"AA9A"
    )
    port map (
      I0 => blk00000001_sig00000e97,
      I1 => blk00000001_sig00000e98,
      I2 => blk00000001_sig00000eac,
      I3 => blk00000001_sig00000eaa,
      O => blk00000001_sig00000e8a
    );
  blk00000001_blk00000c7f : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_sig00000e97,
      I1 => blk00000001_sig00000eaa,
      I2 => blk00000001_sig00000eac,
      O => blk00000001_sig00000e88
    );
  blk00000001_blk00000c7e : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_sig00000e98,
      I1 => blk00000001_sig00000eaa,
      I2 => blk00000001_sig00000eac,
      O => blk00000001_sig00000e89
    );
  blk00000001_blk00000c7d : LUT4
    generic map(
      INIT => X"AA9A"
    )
    port map (
      I0 => blk00000001_sig00000e95,
      I1 => blk00000001_sig00000e96,
      I2 => blk00000001_sig00000eab,
      I3 => blk00000001_sig00000eaa,
      O => blk00000001_sig00000e87
    );
  blk00000001_blk00000c7c : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_sig00000e95,
      I1 => blk00000001_sig00000eaa,
      I2 => blk00000001_sig00000eab,
      O => blk00000001_sig00000e85
    );
  blk00000001_blk00000c7b : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_sig00000e96,
      I1 => blk00000001_sig00000eaa,
      I2 => blk00000001_sig00000eab,
      O => blk00000001_sig00000e86
    );
  blk00000001_blk00000c7a : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => blk00000001_sig00000e9a,
      I1 => blk00000001_sig00000ea1,
      I2 => blk00000001_sig00000ea0,
      O => blk00000001_sig00000e8c
    );
  blk00000001_blk00000c79 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ea1,
      I1 => blk00000001_sig00000ea0,
      O => blk00000001_sig00000e91
    );
  blk00000001_blk00000c78 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000001_sig00000e9a,
      I1 => blk00000001_sig00000ea0,
      I2 => blk00000001_sig00000ea1,
      O => blk00000001_sig00000e8b
    );
  blk00000001_blk00000c77 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_sig00000e9a,
      I1 => blk00000001_sig00000ea0,
      O => blk00000001_sig00000e8d
    );
  blk00000001_blk00000c76 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000e9a,
      I1 => blk00000001_sig00000ea0,
      O => blk00000001_sig00000e90
    );
  blk00000001_blk00000c75 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig000001b0,
      I1 => blk00000001_sig00000e28,
      I2 => blk00000001_sig000001b2,
      I3 => blk00000001_sig00000e2a,
      I4 => blk00000001_sig000001b1,
      I5 => blk00000001_sig00000e29,
      O => blk00000001_sig00000e6d
    );
  blk00000001_blk00000c74 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig000000bb,
      I1 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e0e
    );
  blk00000001_blk00000c73 : LUT3
    generic map(
      INIT => X"40"
    )
    port map (
      I0 => blk00000001_sig00000e1e,
      I1 => blk00000001_sig000000bc,
      I2 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e0c
    );
  blk00000001_blk00000c72 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000e1e,
      I1 => blk00000001_sig000000bc,
      I2 => blk00000001_sig0000008e,
      O => blk00000001_sig00000deb
    );
  blk00000001_blk00000c71 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig000000bb,
      O => blk00000001_sig00000e0b
    );
  blk00000001_blk00000c70 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e22,
      O => blk00000001_sig000001ab
    );
  blk00000001_blk00000c6f : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e21,
      O => blk00000001_sig00000e0a
    );
  blk00000001_blk00000c6e : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig000000bb,
      I1 => blk00000001_sig00000e16,
      O => blk00000001_sig00000dec
    );
  blk00000001_blk00000c6d : LUT4
    generic map(
      INIT => X"EEEF"
    )
    port map (
      I0 => blk00000001_sig00000e1f,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig00000e1d,
      I3 => blk00000001_sig00000e23,
      O => blk00000001_sig00000e09
    );
  blk00000001_blk00000c6c : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000dfb,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000df9
    );
  blk00000001_blk00000c6b : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000dfc,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000dfa
    );
  blk00000001_blk00000c6a : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000dfd,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000df5
    );
  blk00000001_blk00000c69 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000dfe,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000df6
    );
  blk00000001_blk00000c68 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000dff,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000df7
    );
  blk00000001_blk00000c67 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig00000e00,
      I1 => blk00000001_sig00000e11,
      I2 => blk00000001_sig00000e10,
      O => blk00000001_sig00000df8
    );
  blk00000001_blk00000c66 : LUT4
    generic map(
      INIT => X"0E00"
    )
    port map (
      I0 => blk00000001_sig00000e13,
      I1 => blk00000001_sig00000e1f,
      I2 => blk00000001_sig0000008d,
      I3 => blk00000001_sig0000008a,
      O => blk00000001_sig00000dee
    );
  blk00000001_blk00000c65 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig00000e1b,
      I1 => blk00000001_sig00000e1c,
      O => blk00000001_sig00000e05
    );
  blk00000001_blk00000c64 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_sig00000e1b,
      I1 => blk00000001_sig00000e1c,
      O => blk00000001_sig00000e06
    );
  blk00000001_blk00000c63 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_sig00000e1c,
      I1 => blk00000001_sig00000e1b,
      O => blk00000001_sig00000e04
    );
  blk00000001_blk00000c62 : LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000001_sig00000e1b,
      I1 => blk00000001_sig00000e1c,
      O => blk00000001_sig00000e03
    );
  blk00000001_blk00000c61 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig000000bc,
      I1 => blk00000001_sig00000e24,
      I2 => blk00000001_sig00000dea,
      O => blk00000001_sig00000e08
    );
  blk00000001_blk00000c60 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig00000e24,
      I1 => blk00000001_sig00000dea,
      O => blk00000001_sig00000e07
    );
  blk00000001_blk00000c5f : LUT4
    generic map(
      INIT => X"AE00"
    )
    port map (
      I0 => blk00000001_sig000001a8,
      I1 => blk00000001_sig00000e12,
      I2 => blk00000001_sig0000008d,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig00000e0d
    );
  blk00000001_blk00000c5e : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_sig0000008d,
      I1 => blk00000001_sig00000e12,
      O => blk00000001_sig00000ded
    );
  blk00000001_blk00000c5d : LUT6
    generic map(
      INIT => X"56A9A9566A95956A"
    )
    port map (
      I0 => blk00000001_sig00000dfe,
      I1 => blk00000001_sig00000dff,
      I2 => blk00000001_sig00000dfb,
      I3 => blk00000001_sig00000e00,
      I4 => blk00000001_sig00000dfc,
      I5 => blk00000001_sig00000dfd,
      O => blk00000001_sig00000e01
    );
  blk00000001_blk00000c5c : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => blk00000001_sig00000dfd,
      I1 => blk00000001_sig00000dff,
      I2 => blk00000001_sig00000dfb,
      O => blk00000001_sig00000e02
    );
  blk00000001_blk00000c5b : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig00000ddc,
      O => blk00000001_sig000001a5
    );
  blk00000001_blk00000c5a : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig00000ddf,
      I1 => blk00000001_sig0000008e,
      O => blk00000001_sig000001ae
    );
  blk00000001_blk00000c59 : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_sig00000de7,
      I1 => blk00000001_sig00000e1a,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000de0,
      O => blk00000001_sig00000da4
    );
  blk00000001_blk00000c58 : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_sig00000de7,
      I1 => blk00000001_sig00000e19,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000de0,
      O => blk00000001_sig00000da3
    );
  blk00000001_blk00000c57 : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_sig00000de7,
      I1 => blk00000001_sig00000e18,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000de0,
      O => blk00000001_sig00000da2
    );
  blk00000001_blk00000c56 : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_sig00000de7,
      I1 => blk00000001_sig00000e17,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig00000de0,
      O => blk00000001_sig00000da1
    );
  blk00000001_blk00000c55 : LUT3
    generic map(
      INIT => X"4E"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      O => blk00000001_sig00000cd1
    );
  blk00000001_blk00000c54 : LUT3
    generic map(
      INIT => X"1B"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      O => blk00000001_sig00000cd0
    );
  blk00000001_blk00000c53 : LUT3
    generic map(
      INIT => X"A9"
    )
    port map (
      I0 => blk00000001_sig000001b5,
      I1 => blk00000001_sig000001ac,
      I2 => blk00000001_sig000001b6,
      O => blk00000001_sig00000ccf
    );
  blk00000001_blk00000c52 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_sig000001b5,
      I1 => blk00000001_sig000001ac,
      I2 => blk00000001_sig000001b6,
      O => blk00000001_sig00000cce
    );
  blk00000001_blk00000c51 : LUT4
    generic map(
      INIT => X"78D8"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      I3 => blk00000001_sig000001e0,
      O => blk00000001_sig00000cd2
    );
  blk00000001_blk00000c50 : LUT4
    generic map(
      INIT => X"8D87"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      I3 => blk00000001_sig000001e0,
      O => blk00000001_sig00000ccd
    );
  blk00000001_blk00000c4f : LUT4
    generic map(
      INIT => X"D272"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      I3 => blk00000001_sig000001e0,
      O => blk00000001_sig00000ccb
    );
  blk00000001_blk00000c4e : LUT4
    generic map(
      INIT => X"272D"
    )
    port map (
      I0 => blk00000001_sig000001ac,
      I1 => blk00000001_sig000001b6,
      I2 => blk00000001_sig000001b5,
      I3 => blk00000001_sig000001e0,
      O => blk00000001_sig00000ccc
    );
  blk00000001_blk00000c4d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005cf,
      I2 => blk00000001_sig0000060b,
      O => blk00000001_sig00000c1f
    );
  blk00000001_blk00000c4c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005ce,
      I2 => blk00000001_sig0000060a,
      O => blk00000001_sig00000c1e
    );
  blk00000001_blk00000c4b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005cd,
      I2 => blk00000001_sig00000609,
      O => blk00000001_sig00000c1d
    );
  blk00000001_blk00000c4a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005cc,
      I2 => blk00000001_sig00000608,
      O => blk00000001_sig00000c1c
    );
  blk00000001_blk00000c49 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005cb,
      I2 => blk00000001_sig00000607,
      O => blk00000001_sig00000c1b
    );
  blk00000001_blk00000c48 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005ca,
      I2 => blk00000001_sig00000606,
      O => blk00000001_sig00000c1a
    );
  blk00000001_blk00000c47 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c9,
      I2 => blk00000001_sig00000605,
      O => blk00000001_sig00000c19
    );
  blk00000001_blk00000c46 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c8,
      I2 => blk00000001_sig00000604,
      O => blk00000001_sig00000c18
    );
  blk00000001_blk00000c45 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d9,
      I2 => blk00000001_sig00000615,
      O => blk00000001_sig00000c29
    );
  blk00000001_blk00000c44 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d8,
      I2 => blk00000001_sig00000614,
      O => blk00000001_sig00000c28
    );
  blk00000001_blk00000c43 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d7,
      I2 => blk00000001_sig00000613,
      O => blk00000001_sig00000c27
    );
  blk00000001_blk00000c42 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d6,
      I2 => blk00000001_sig00000612,
      O => blk00000001_sig00000c26
    );
  blk00000001_blk00000c41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d5,
      I2 => blk00000001_sig00000611,
      O => blk00000001_sig00000c25
    );
  blk00000001_blk00000c40 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d4,
      I2 => blk00000001_sig00000610,
      O => blk00000001_sig00000c24
    );
  blk00000001_blk00000c3f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d3,
      I2 => blk00000001_sig0000060f,
      O => blk00000001_sig00000c23
    );
  blk00000001_blk00000c3e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d2,
      I2 => blk00000001_sig0000060e,
      O => blk00000001_sig00000c22
    );
  blk00000001_blk00000c3d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d1,
      I2 => blk00000001_sig0000060d,
      O => blk00000001_sig00000c21
    );
  blk00000001_blk00000c3c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005d0,
      I2 => blk00000001_sig0000060c,
      O => blk00000001_sig00000c20
    );
  blk00000001_blk00000c3b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c7,
      I2 => blk00000001_sig00000603,
      O => blk00000001_sig00000c17
    );
  blk00000001_blk00000c3a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c6,
      I2 => blk00000001_sig00000602,
      O => blk00000001_sig00000c16
    );
  blk00000001_blk00000c39 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005bb,
      I2 => blk00000001_sig000005cf,
      O => blk00000001_sig00000c0b
    );
  blk00000001_blk00000c38 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005ba,
      I2 => blk00000001_sig000005ce,
      O => blk00000001_sig00000c0a
    );
  blk00000001_blk00000c37 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b9,
      I2 => blk00000001_sig000005cd,
      O => blk00000001_sig00000c09
    );
  blk00000001_blk00000c36 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b8,
      I2 => blk00000001_sig000005cc,
      O => blk00000001_sig00000c08
    );
  blk00000001_blk00000c35 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b7,
      I2 => blk00000001_sig000005cb,
      O => blk00000001_sig00000c07
    );
  blk00000001_blk00000c34 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b6,
      I2 => blk00000001_sig000005ca,
      O => blk00000001_sig00000c06
    );
  blk00000001_blk00000c33 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b5,
      I2 => blk00000001_sig000005c9,
      O => blk00000001_sig00000c05
    );
  blk00000001_blk00000c32 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b4,
      I2 => blk00000001_sig000005c8,
      O => blk00000001_sig00000c04
    );
  blk00000001_blk00000c31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c5,
      I2 => blk00000001_sig000005d9,
      O => blk00000001_sig00000c15
    );
  blk00000001_blk00000c30 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c4,
      I2 => blk00000001_sig000005d8,
      O => blk00000001_sig00000c14
    );
  blk00000001_blk00000c2f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c3,
      I2 => blk00000001_sig000005d7,
      O => blk00000001_sig00000c13
    );
  blk00000001_blk00000c2e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c2,
      I2 => blk00000001_sig000005d6,
      O => blk00000001_sig00000c12
    );
  blk00000001_blk00000c2d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c1,
      I2 => blk00000001_sig000005d5,
      O => blk00000001_sig00000c11
    );
  blk00000001_blk00000c2c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005c0,
      I2 => blk00000001_sig000005d4,
      O => blk00000001_sig00000c10
    );
  blk00000001_blk00000c2b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005bf,
      I2 => blk00000001_sig000005d3,
      O => blk00000001_sig00000c0f
    );
  blk00000001_blk00000c2a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005be,
      I2 => blk00000001_sig000005d2,
      O => blk00000001_sig00000c0e
    );
  blk00000001_blk00000c29 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005bd,
      I2 => blk00000001_sig000005d1,
      O => blk00000001_sig00000c0d
    );
  blk00000001_blk00000c28 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005bc,
      I2 => blk00000001_sig000005d0,
      O => blk00000001_sig00000c0c
    );
  blk00000001_blk00000c27 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b3,
      I2 => blk00000001_sig000005c7,
      O => blk00000001_sig00000c03
    );
  blk00000001_blk00000c26 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig00000ba0,
      I1 => blk00000001_sig000005b2,
      I2 => blk00000001_sig000005c6,
      O => blk00000001_sig00000c02
    );
  blk00000001_blk00000c25 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig0000008e,
      I1 => blk00000001_sig0000008b,
      O => blk00000001_sig000002e3
    );
  blk00000001_blk00000c24 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig000001e0,
      I1 => blk00000001_sig000002e1,
      O => blk00000001_sig000001d9
    );
  blk00000001_blk00000c23 : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => NlwRenamedSig_OI_s_axis_data_tready,
      I1 => aclken,
      I2 => blk00000001_sig000000f8,
      I3 => s_axis_data_tvalid,
      O => blk00000001_sig00000180
    );
  blk00000001_blk00000c22 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_s_axis_data_tready,
      I2 => blk00000001_sig00000182,
      O => blk00000001_sig0000017f
    );
  blk00000001_blk00000c21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000167,
      I2 => blk00000001_sig00000144,
      O => blk00000001_sig00000121
    );
  blk00000001_blk00000c20 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000166,
      I2 => blk00000001_sig00000143,
      O => blk00000001_sig00000120
    );
  blk00000001_blk00000c1f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000165,
      I2 => blk00000001_sig00000142,
      O => blk00000001_sig0000011f
    );
  blk00000001_blk00000c1e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000164,
      I2 => blk00000001_sig00000141,
      O => blk00000001_sig0000011e
    );
  blk00000001_blk00000c1d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000163,
      I2 => blk00000001_sig00000140,
      O => blk00000001_sig0000011d
    );
  blk00000001_blk00000c1c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000162,
      I2 => blk00000001_sig0000013f,
      O => blk00000001_sig0000011c
    );
  blk00000001_blk00000c1b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000017e,
      I2 => blk00000001_sig0000015b,
      O => blk00000001_sig00000138
    );
  blk00000001_blk00000c1a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000017d,
      I2 => blk00000001_sig0000015a,
      O => blk00000001_sig00000137
    );
  blk00000001_blk00000c19 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000017c,
      I2 => blk00000001_sig00000159,
      O => blk00000001_sig00000136
    );
  blk00000001_blk00000c18 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000161,
      I2 => blk00000001_sig0000013e,
      O => blk00000001_sig0000011b
    );
  blk00000001_blk00000c17 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000017b,
      I2 => blk00000001_sig00000158,
      O => blk00000001_sig00000135
    );
  blk00000001_blk00000c16 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000017a,
      I2 => blk00000001_sig00000157,
      O => blk00000001_sig00000134
    );
  blk00000001_blk00000c15 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000179,
      I2 => blk00000001_sig00000156,
      O => blk00000001_sig00000133
    );
  blk00000001_blk00000c14 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000178,
      I2 => blk00000001_sig00000155,
      O => blk00000001_sig00000132
    );
  blk00000001_blk00000c13 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000177,
      I2 => blk00000001_sig00000154,
      O => blk00000001_sig00000131
    );
  blk00000001_blk00000c12 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000176,
      I2 => blk00000001_sig00000153,
      O => blk00000001_sig00000130
    );
  blk00000001_blk00000c11 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000175,
      I2 => blk00000001_sig00000152,
      O => blk00000001_sig0000012f
    );
  blk00000001_blk00000c10 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000174,
      I2 => blk00000001_sig00000151,
      O => blk00000001_sig0000012e
    );
  blk00000001_blk00000c0f : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000173,
      I2 => blk00000001_sig00000150,
      O => blk00000001_sig0000012d
    );
  blk00000001_blk00000c0e : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000172,
      I2 => blk00000001_sig0000014f,
      O => blk00000001_sig0000012c
    );
  blk00000001_blk00000c0d : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000160,
      I2 => blk00000001_sig0000013d,
      O => blk00000001_sig0000011a
    );
  blk00000001_blk00000c0c : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000171,
      I2 => blk00000001_sig0000014e,
      O => blk00000001_sig0000012b
    );
  blk00000001_blk00000c0b : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000170,
      I2 => blk00000001_sig0000014d,
      O => blk00000001_sig0000012a
    );
  blk00000001_blk00000c0a : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016f,
      I2 => blk00000001_sig0000014c,
      O => blk00000001_sig00000129
    );
  blk00000001_blk00000c09 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016e,
      I2 => blk00000001_sig0000014b,
      O => blk00000001_sig00000128
    );
  blk00000001_blk00000c08 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016d,
      I2 => blk00000001_sig0000014a,
      O => blk00000001_sig00000127
    );
  blk00000001_blk00000c07 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016c,
      I2 => blk00000001_sig00000149,
      O => blk00000001_sig00000126
    );
  blk00000001_blk00000c06 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016b,
      I2 => blk00000001_sig00000148,
      O => blk00000001_sig00000125
    );
  blk00000001_blk00000c05 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000016a,
      I2 => blk00000001_sig00000147,
      O => blk00000001_sig00000124
    );
  blk00000001_blk00000c04 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000169,
      I2 => blk00000001_sig00000146,
      O => blk00000001_sig00000123
    );
  blk00000001_blk00000c03 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig00000168,
      I2 => blk00000001_sig00000145,
      O => blk00000001_sig00000122
    );
  blk00000001_blk00000c02 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000015f,
      I2 => blk00000001_sig0000013c,
      O => blk00000001_sig00000119
    );
  blk00000001_blk00000c01 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig0000013a,
      I1 => blk00000001_sig0000015e,
      I2 => blk00000001_sig0000013b,
      O => blk00000001_sig00000118
    );
  blk00000001_blk00000c00 : LUT4
    generic map(
      INIT => X"FA32"
    )
    port map (
      I0 => blk00000001_sig0000015c,
      I1 => blk00000001_sig00000101,
      I2 => blk00000001_sig0000013a,
      I3 => blk00000001_sig000000dc,
      O => blk00000001_sig00000116
    );
  blk00000001_blk00000bff : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => NlwRenamedSig_OI_s_axis_config_tready,
      I1 => aclken,
      I2 => blk00000001_sig000000f8,
      I3 => s_axis_config_tvalid,
      O => blk00000001_sig0000010c
    );
  blk00000001_blk00000bfe : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_s_axis_config_tready,
      I2 => blk00000001_sig0000010e,
      O => blk00000001_sig0000010b
    );
  blk00000001_blk00000bfd : LUT6
    generic map(
      INIT => X"EAEAC0C0FFEAFFC0"
    )
    port map (
      I0 => blk00000001_sig000000e2,
      I1 => blk00000001_sig000000e0,
      I2 => blk00000001_sig000000bd,
      I3 => blk00000001_sig000000e1,
      I4 => blk00000001_sig00000101,
      I5 => blk00000001_sig000000bb,
      O => blk00000001_sig0000008a
    );
  blk00000001_blk00000bfc : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_sig000000be,
      I1 => blk00000001_sig000000de,
      O => blk00000001_sig000000d3
    );
  blk00000001_blk00000bfb : LUT3
    generic map(
      INIT => X"F2"
    )
    port map (
      I0 => blk00000001_sig000000e2,
      I1 => blk00000001_sig00000101,
      I2 => blk00000001_sig000000e3,
      O => blk00000001_sig000000d0
    );
  blk00000001_blk00000bfa : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig0000010a,
      I2 => blk00000001_sig000000ea,
      O => blk00000001_sig00000078
    );
  blk00000001_blk00000bf9 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000109,
      I2 => blk00000001_sig000000e9,
      O => blk00000001_sig00000079
    );
  blk00000001_blk00000bf8 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000108,
      I2 => blk00000001_sig000000e8,
      O => blk00000001_sig0000007a
    );
  blk00000001_blk00000bf7 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000107,
      I2 => blk00000001_sig000000e7,
      O => blk00000001_sig0000007b
    );
  blk00000001_blk00000bf6 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000106,
      I2 => blk00000001_sig000000e6,
      O => blk00000001_sig0000007c
    );
  blk00000001_blk00000bf5 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000105,
      I2 => blk00000001_sig000000e5,
      O => blk00000001_sig0000007d
    );
  blk00000001_blk00000bf4 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => blk00000001_sig000000e3,
      I1 => blk00000001_sig00000104,
      I2 => blk00000001_sig000000e4,
      O => blk00000001_sig0000008c
    );
  blk00000001_blk00000bf3 : LUT6
    generic map(
      INIT => X"7FFFFFFFFFFFFFFF"
    )
    port map (
      I0 => blk00000001_sig00000092,
      I1 => blk00000001_sig00000091,
      I2 => blk00000001_sig00000090,
      I3 => blk00000001_sig0000008f,
      I4 => blk00000001_sig00000094,
      I5 => blk00000001_sig00000093,
      O => blk00000001_sig000000c5
    );
  blk00000001_blk00000bf2 : LUT5
    generic map(
      INIT => X"AA00EAC0"
    )
    port map (
      I0 => blk00000001_sig000000de,
      I1 => blk00000001_sig000000df,
      I2 => blk00000001_sig000000f3,
      I3 => blk00000001_sig000000be,
      I4 => blk00000001_sig000000c5,
      O => blk00000001_sig000000d4
    );
  blk00000001_blk00000bf1 : LUT5
    generic map(
      INIT => X"222222F2"
    )
    port map (
      I0 => blk00000001_sig000000e0,
      I1 => blk00000001_sig000000bd,
      I2 => blk00000001_sig000000df,
      I3 => blk00000001_sig000000f3,
      I4 => blk00000001_sig000000c5,
      O => blk00000001_sig000000ce
    );
  blk00000001_blk00000bf0 : LUT5
    generic map(
      INIT => X"00000001"
    )
    port map (
      I0 => blk00000001_sig000000ee,
      I1 => blk00000001_sig000000ef,
      I2 => blk00000001_sig000000f0,
      I3 => blk00000001_sig000000f1,
      I4 => blk00000001_sig000000f2,
      O => blk00000001_sig000000c4
    );
  blk00000001_blk00000bef : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => blk00000001_sig000000f3,
      I1 => blk00000001_sig00000fcb,
      O => blk00000001_sig000000c3
    );
  blk00000001_blk00000bee : LUT3
    generic map(
      INIT => X"20"
    )
    port map (
      I0 => blk00000001_sig000000be,
      I1 => blk00000001_sig000000f8,
      I2 => blk00000001_sig0000008e,
      O => blk00000001_sig000000da
    );
  blk00000001_blk00000bed : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig000000be,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000c4,
      O => blk00000001_sig000000db
    );
  blk00000001_blk00000bec : LUT6
    generic map(
      INIT => X"008800A800000000"
    )
    port map (
      I0 => blk00000001_sig000000e0,
      I1 => blk00000001_sig000000bd,
      I2 => blk00000001_sig000000e1,
      I3 => blk00000001_sig00000101,
      I4 => blk00000001_sig000000bb,
      I5 => blk00000001_sig0000008e,
      O => blk00000001_sig000000d6
    );
  blk00000001_blk00000beb : LUT5
    generic map(
      INIT => X"73005000"
    )
    port map (
      I0 => blk00000001_sig000000f4,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000be,
      I3 => blk00000001_sig0000008e,
      I4 => blk00000001_sig000000c4,
      O => blk00000001_sig000000d7
    );
  blk00000001_blk00000bea : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig000000df,
      I1 => blk00000001_sig000000c5,
      O => blk00000001_sig000000c1
    );
  blk00000001_blk00000be9 : LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      I0 => blk00000001_sig000000f3,
      I1 => blk00000001_sig000000bb,
      I2 => blk00000001_sig000000f8,
      I3 => blk00000001_sig00000fcb,
      O => blk00000001_sig000000dc
    );
  blk00000001_blk00000be8 : LUT6
    generic map(
      INIT => X"CCECCCECCCECCCCC"
    )
    port map (
      I0 => blk00000001_sig000000f5,
      I1 => blk00000001_sig000000dd,
      I2 => blk00000001_sig000000e1,
      I3 => blk00000001_sig000000f3,
      I4 => blk00000001_sig000000bb,
      I5 => blk00000001_sig000000c1,
      O => blk00000001_sig000000d1
    );
  blk00000001_blk00000be7 : LUT3
    generic map(
      INIT => X"20"
    )
    port map (
      I0 => blk00000001_sig000000fa,
      I1 => blk00000001_sig00000100,
      I2 => blk00000001_sig0000008e,
      O => blk00000001_sig000000d8
    );
  blk00000001_blk00000be6 : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => blk00000001_sig000000eb,
      I1 => blk00000001_sig000000fa,
      I2 => blk00000001_sig00000100,
      I3 => blk00000001_sig0000008e,
      O => blk00000001_sig000000cb
    );
  blk00000001_blk00000be5 : LUT5
    generic map(
      INIT => X"DFFF8AAA"
    )
    port map (
      I0 => blk00000001_sig000000eb,
      I1 => blk00000001_sig00000100,
      I2 => blk00000001_sig0000008e,
      I3 => blk00000001_sig000000fa,
      I4 => blk00000001_sig000000db,
      O => blk00000001_sig000000d2
    );
  blk00000001_blk00000be4 : LUT5
    generic map(
      INIT => X"AAAAAAA9"
    )
    port map (
      I0 => blk00000001_sig000000f1,
      I1 => blk00000001_sig000000c6,
      I2 => blk00000001_sig000000ee,
      I3 => blk00000001_sig000000ef,
      I4 => blk00000001_sig000000f0,
      O => blk00000001_sig000000ca
    );
  blk00000001_blk00000be3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f59,
      Q => blk00000001_sig000008d0
    );
  blk00000001_blk00000be2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5a,
      Q => blk00000001_sig000008d1
    );
  blk00000001_blk00000be1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5b,
      Q => blk00000001_sig000008d2
    );
  blk00000001_blk00000be0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5c,
      Q => blk00000001_sig000008d3
    );
  blk00000001_blk00000bdf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5d,
      Q => blk00000001_sig000008d4
    );
  blk00000001_blk00000bde : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5e,
      Q => blk00000001_sig000008d5
    );
  blk00000001_blk00000bdd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f5f,
      Q => blk00000001_sig000008d6
    );
  blk00000001_blk00000bdc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f60,
      Q => blk00000001_sig000008d7
    );
  blk00000001_blk00000bdb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f61,
      Q => blk00000001_sig000008d8
    );
  blk00000001_blk00000bda : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f62,
      Q => blk00000001_sig000008d9
    );
  blk00000001_blk00000bd9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f63,
      Q => blk00000001_sig000008da
    );
  blk00000001_blk00000bd8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f64,
      Q => blk00000001_sig000008db
    );
  blk00000001_blk00000bd7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f65,
      Q => blk00000001_sig000008dc
    );
  blk00000001_blk00000bd6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f66,
      Q => blk00000001_sig000008dd
    );
  blk00000001_blk00000bd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f67,
      Q => blk00000001_sig000008de
    );
  blk00000001_blk00000bd4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f68,
      Q => blk00000001_sig000008df
    );
  blk00000001_blk00000bd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f69,
      Q => blk00000001_sig000008e0
    );
  blk00000001_blk00000bd2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f48,
      Q => blk00000001_sig000008e1
    );
  blk00000001_blk00000bd1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f49,
      Q => blk00000001_sig000008e2
    );
  blk00000001_blk00000bd0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4a,
      Q => blk00000001_sig000008e3
    );
  blk00000001_blk00000bcf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4b,
      Q => blk00000001_sig000008e4
    );
  blk00000001_blk00000bce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4c,
      Q => blk00000001_sig000008e5
    );
  blk00000001_blk00000bcd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4d,
      Q => blk00000001_sig000008e6
    );
  blk00000001_blk00000bcc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4e,
      Q => blk00000001_sig000008e7
    );
  blk00000001_blk00000bcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f4f,
      Q => blk00000001_sig000008e8
    );
  blk00000001_blk00000bca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f50,
      Q => blk00000001_sig000008e9
    );
  blk00000001_blk00000bc9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f51,
      Q => blk00000001_sig000008ea
    );
  blk00000001_blk00000bc8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f52,
      Q => blk00000001_sig000008eb
    );
  blk00000001_blk00000bc7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f53,
      Q => blk00000001_sig000008ec
    );
  blk00000001_blk00000bc6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f54,
      Q => blk00000001_sig000008ed
    );
  blk00000001_blk00000bc5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f55,
      Q => blk00000001_sig000008ee
    );
  blk00000001_blk00000bc4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f56,
      Q => blk00000001_sig000008ef
    );
  blk00000001_blk00000bc3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f57,
      Q => blk00000001_sig000008f0
    );
  blk00000001_blk00000bc2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f58,
      Q => blk00000001_sig000008f1
    );
  blk00000001_blk00000bc1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f37,
      Q => blk00000001_sig0000085b
    );
  blk00000001_blk00000bc0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f38,
      Q => blk00000001_sig0000085c
    );
  blk00000001_blk00000bbf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f39,
      Q => blk00000001_sig0000085d
    );
  blk00000001_blk00000bbe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3a,
      Q => blk00000001_sig0000085e
    );
  blk00000001_blk00000bbd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3b,
      Q => blk00000001_sig0000085f
    );
  blk00000001_blk00000bbc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3c,
      Q => blk00000001_sig00000860
    );
  blk00000001_blk00000bbb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3d,
      Q => blk00000001_sig00000861
    );
  blk00000001_blk00000bba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3e,
      Q => blk00000001_sig00000862
    );
  blk00000001_blk00000bb9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f3f,
      Q => blk00000001_sig00000863
    );
  blk00000001_blk00000bb8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f40,
      Q => blk00000001_sig00000864
    );
  blk00000001_blk00000bb7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f41,
      Q => blk00000001_sig00000865
    );
  blk00000001_blk00000bb6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f42,
      Q => blk00000001_sig00000866
    );
  blk00000001_blk00000bb5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f43,
      Q => blk00000001_sig00000867
    );
  blk00000001_blk00000bb4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f44,
      Q => blk00000001_sig00000868
    );
  blk00000001_blk00000bb3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f45,
      Q => blk00000001_sig00000869
    );
  blk00000001_blk00000bb2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f46,
      Q => blk00000001_sig0000086a
    );
  blk00000001_blk00000bb1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f47,
      Q => blk00000001_sig0000086b
    );
  blk00000001_blk00000bb0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f26,
      Q => blk00000001_sig0000086c
    );
  blk00000001_blk00000baf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f27,
      Q => blk00000001_sig0000086d
    );
  blk00000001_blk00000bae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f28,
      Q => blk00000001_sig0000086e
    );
  blk00000001_blk00000bad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f29,
      Q => blk00000001_sig0000086f
    );
  blk00000001_blk00000bac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2a,
      Q => blk00000001_sig00000870
    );
  blk00000001_blk00000bab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2b,
      Q => blk00000001_sig00000871
    );
  blk00000001_blk00000baa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2c,
      Q => blk00000001_sig00000872
    );
  blk00000001_blk00000ba9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2d,
      Q => blk00000001_sig00000873
    );
  blk00000001_blk00000ba8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2e,
      Q => blk00000001_sig00000874
    );
  blk00000001_blk00000ba7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f2f,
      Q => blk00000001_sig00000875
    );
  blk00000001_blk00000ba6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f30,
      Q => blk00000001_sig00000876
    );
  blk00000001_blk00000ba5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f31,
      Q => blk00000001_sig00000877
    );
  blk00000001_blk00000ba4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f32,
      Q => blk00000001_sig00000878
    );
  blk00000001_blk00000ba3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f33,
      Q => blk00000001_sig00000879
    );
  blk00000001_blk00000ba2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f34,
      Q => blk00000001_sig0000087a
    );
  blk00000001_blk00000ba1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f35,
      Q => blk00000001_sig0000087b
    );
  blk00000001_blk00000ba0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f36,
      Q => blk00000001_sig0000087c
    );
  blk00000001_blk00000b9f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f15,
      Q => blk00000001_sig000007e8
    );
  blk00000001_blk00000b9e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f16,
      Q => blk00000001_sig000007e9
    );
  blk00000001_blk00000b9d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f17,
      Q => blk00000001_sig000007ea
    );
  blk00000001_blk00000b9c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f18,
      Q => blk00000001_sig000007eb
    );
  blk00000001_blk00000b9b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f19,
      Q => blk00000001_sig000007ec
    );
  blk00000001_blk00000b9a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1a,
      Q => blk00000001_sig000007ed
    );
  blk00000001_blk00000b99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1b,
      Q => blk00000001_sig000007ee
    );
  blk00000001_blk00000b98 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1c,
      Q => blk00000001_sig000007ef
    );
  blk00000001_blk00000b97 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1d,
      Q => blk00000001_sig000007f0
    );
  blk00000001_blk00000b96 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1e,
      Q => blk00000001_sig000007f1
    );
  blk00000001_blk00000b95 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f1f,
      Q => blk00000001_sig000007f2
    );
  blk00000001_blk00000b94 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f20,
      Q => blk00000001_sig000007f3
    );
  blk00000001_blk00000b93 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f21,
      Q => blk00000001_sig000007f4
    );
  blk00000001_blk00000b92 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f22,
      Q => blk00000001_sig000007f5
    );
  blk00000001_blk00000b91 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f23,
      Q => blk00000001_sig000007f6
    );
  blk00000001_blk00000b90 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f24,
      Q => blk00000001_sig000007f7
    );
  blk00000001_blk00000b8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f25,
      Q => blk00000001_sig000007f8
    );
  blk00000001_blk00000b8e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f04,
      Q => blk00000001_sig000007f9
    );
  blk00000001_blk00000b8d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f05,
      Q => blk00000001_sig000007fa
    );
  blk00000001_blk00000b8c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f06,
      Q => blk00000001_sig000007fb
    );
  blk00000001_blk00000b8b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f07,
      Q => blk00000001_sig000007fc
    );
  blk00000001_blk00000b8a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f08,
      Q => blk00000001_sig000007fd
    );
  blk00000001_blk00000b89 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f09,
      Q => blk00000001_sig000007fe
    );
  blk00000001_blk00000b88 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0a,
      Q => blk00000001_sig000007ff
    );
  blk00000001_blk00000b87 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0b,
      Q => blk00000001_sig00000800
    );
  blk00000001_blk00000b86 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0c,
      Q => blk00000001_sig00000801
    );
  blk00000001_blk00000b85 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0d,
      Q => blk00000001_sig00000802
    );
  blk00000001_blk00000b84 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0e,
      Q => blk00000001_sig00000803
    );
  blk00000001_blk00000b83 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f0f,
      Q => blk00000001_sig00000804
    );
  blk00000001_blk00000b82 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f10,
      Q => blk00000001_sig00000805
    );
  blk00000001_blk00000b81 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f11,
      Q => blk00000001_sig00000806
    );
  blk00000001_blk00000b80 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f12,
      Q => blk00000001_sig00000807
    );
  blk00000001_blk00000b7f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f13,
      Q => blk00000001_sig00000808
    );
  blk00000001_blk00000b7e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f14,
      Q => blk00000001_sig00000809
    );
  blk00000001_blk00000b3b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f03,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000eff
    );
  blk00000001_blk00000b3a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f02,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000efe
    );
  blk00000001_blk00000b39 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f01,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000efd
    );
  blk00000001_blk00000b38 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000f00,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000efc
    );
  blk00000001_blk00000b37 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000de4,
      I2 => blk00000001_sig00000de6,
      I3 => blk00000001_sig00000de1,
      I4 => blk00000001_sig00000de2,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000f03
    );
  blk00000001_blk00000b36 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000de3,
      I2 => blk00000001_sig00000de5,
      I3 => blk00000001_sig00000de1,
      I4 => blk00000001_sig00000de2,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000f02
    );
  blk00000001_blk00000b35 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000de4,
      I3 => blk00000001_sig00000de1,
      I4 => blk00000001_sig00000de2,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000f01
    );
  blk00000001_blk00000b34 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000de3,
      I3 => blk00000001_sig00000de1,
      I4 => blk00000001_sig00000de2,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000f00
    );
  blk00000001_blk00000b33 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef5,
      Q => blk00000001_sig00000dc5
    );
  blk00000001_blk00000b32 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef4,
      Q => blk00000001_sig00000dc6
    );
  blk00000001_blk00000b31 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef3,
      Q => blk00000001_sig00000dc7
    );
  blk00000001_blk00000b30 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef2,
      Q => blk00000001_sig00000dc8
    );
  blk00000001_blk00000b2f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dc9
    );
  blk00000001_blk00000b2e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dc0
    );
  blk00000001_blk00000b2d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef5,
      Q => blk00000001_sig00000dc1
    );
  blk00000001_blk00000b2c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef4,
      Q => blk00000001_sig00000dc2
    );
  blk00000001_blk00000b2b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef3,
      Q => blk00000001_sig00000dc3
    );
  blk00000001_blk00000b2a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef2,
      Q => blk00000001_sig00000dc4
    );
  blk00000001_blk00000b29 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000efb,
      Q => blk00000001_sig000001a6
    );
  blk00000001_blk00000b28 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000efa,
      Q => blk00000001_sig00000dbf
    );
  blk00000001_blk00000b27 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef9,
      Q => blk00000001_sig00000dbe
    );
  blk00000001_blk00000b26 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef8,
      Q => blk00000001_sig00000dbd
    );
  blk00000001_blk00000b25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef7,
      Q => blk00000001_sig00000dbc
    );
  blk00000001_blk00000b24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef6,
      Q => blk00000001_sig00000dbb
    );
  blk00000001_blk00000b23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef1,
      Q => blk00000001_sig00000eea
    );
  blk00000001_blk00000b22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ef0,
      Q => blk00000001_sig00000eeb
    );
  blk00000001_blk00000b21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eef,
      Q => blk00000001_sig00000eec
    );
  blk00000001_blk00000b20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eee,
      Q => blk00000001_sig00000eed
    );
  blk00000001_blk00000b1f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dfd,
      I1 => blk00000001_sig00000dfd,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ef1
    );
  blk00000001_blk00000b1e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dfe,
      I1 => blk00000001_sig00000dfe,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ef0
    );
  blk00000001_blk00000b1d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dff,
      I1 => blk00000001_sig00000dff,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000eef
    );
  blk00000001_blk00000b1c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e00,
      I1 => blk00000001_sig00000e00,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000eee
    );
  blk00000001_blk00000b1b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dfb,
      I1 => blk00000001_sig00000dfb,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000b1b_O_UNCONNECTED
    );
  blk00000001_blk00000b1a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dfc,
      I1 => blk00000001_sig00000dfc,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000b1a_O_UNCONNECTED
    );
  blk00000001_blk00000b19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eea,
      Q => blk00000001_sig00000dca
    );
  blk00000001_blk00000b18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eeb,
      Q => blk00000001_sig00000dcb
    );
  blk00000001_blk00000b17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eec,
      Q => blk00000001_sig00000dcc
    );
  blk00000001_blk00000b16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eed,
      Q => blk00000001_sig00000dcd
    );
  blk00000001_blk00000b15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee9,
      Q => blk00000001_sig00000dce
    );
  blk00000001_blk00000b14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee8,
      Q => blk00000001_sig00000dcf
    );
  blk00000001_blk00000b13 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000ea7,
      I1 => blk00000001_sig00000ea1,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ee9
    );
  blk00000001_blk00000b12 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e92,
      I1 => blk00000001_sig00000e91,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ee8
    );
  blk00000001_blk00000b11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c2
    );
  blk00000001_blk00000b10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c4
    );
  blk00000001_blk00000b0f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd0,
      I1 => blk00000001_sig00000dca,
      I2 => blk00000001_sig00000dde,
      O => NLW_blk00000001_blk00000b0f_O_UNCONNECTED
    );
  blk00000001_blk00000b0e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd1,
      I1 => blk00000001_sig00000dcb,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ee7
    );
  blk00000001_blk00000b0d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd2,
      I1 => blk00000001_sig00000dcc,
      I2 => blk00000001_sig00000dde,
      O => NLW_blk00000001_blk00000b0d_O_UNCONNECTED
    );
  blk00000001_blk00000b0c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd3,
      I1 => blk00000001_sig00000dcd,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ee6
    );
  blk00000001_blk00000b0b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001d1
    );
  blk00000001_blk00000b0a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001d2
    );
  blk00000001_blk00000b09 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001d3
    );
  blk00000001_blk00000b08 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001d4
    );
  blk00000001_blk00000b07 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db3,
      I1 => blk00000001_sig00000db7,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ee5
    );
  blk00000001_blk00000b06 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db4,
      I1 => blk00000001_sig00000db8,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ee4
    );
  blk00000001_blk00000b05 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db5,
      I1 => blk00000001_sig00000db9,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ee3
    );
  blk00000001_blk00000b04 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db6,
      I1 => blk00000001_sig00000dba,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ee2
    );
  blk00000001_blk00000b03 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001be
    );
  blk00000001_blk00000b02 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ee0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c0
    );
  blk00000001_blk00000b01 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd9,
      I1 => blk00000001_sig00000dca,
      I2 => blk00000001_sig00000dde,
      O => NLW_blk00000001_blk00000b01_O_UNCONNECTED
    );
  blk00000001_blk00000b00 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd4,
      I1 => blk00000001_sig00000dcb,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ee1
    );
  blk00000001_blk00000aff : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd5,
      I1 => blk00000001_sig00000dcc,
      I2 => blk00000001_sig00000dde,
      O => NLW_blk00000001_blk00000aff_O_UNCONNECTED
    );
  blk00000001_blk00000afe : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd6,
      I1 => blk00000001_sig00000dcd,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ee0
    );
  blk00000001_blk00000afd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000edf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001cd
    );
  blk00000001_blk00000afc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ede,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001ce
    );
  blk00000001_blk00000afb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000edd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001cf
    );
  blk00000001_blk00000afa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000edc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001d0
    );
  blk00000001_blk00000af9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000daf,
      I1 => blk00000001_sig00000db7,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000edf
    );
  blk00000001_blk00000af8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db0,
      I1 => blk00000001_sig00000db8,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ede
    );
  blk00000001_blk00000af7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db1,
      I1 => blk00000001_sig00000db9,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000edd
    );
  blk00000001_blk00000af6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000db2,
      I1 => blk00000001_sig00000dba,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000edc
    );
  blk00000001_blk00000af5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000edb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c1
    );
  blk00000001_blk00000af4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eda,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001bc
    );
  blk00000001_blk00000af3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c3
    );
  blk00000001_blk00000af2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001bd
    );
  blk00000001_blk00000af1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd0,
      I1 => blk00000001_sig00000dca,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000edb
    );
  blk00000001_blk00000af0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd7,
      I1 => blk00000001_sig00000dcb,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000eda
    );
  blk00000001_blk00000aef : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd2,
      I1 => blk00000001_sig00000dcc,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed9
    );
  blk00000001_blk00000aee : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd8,
      I1 => blk00000001_sig00000dcd,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed8
    );
  blk00000001_blk00000aed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c9
    );
  blk00000001_blk00000aec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001ca
    );
  blk00000001_blk00000aeb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001cb
    );
  blk00000001_blk00000aea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001cc
    );
  blk00000001_blk00000ae9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dab,
      I1 => blk00000001_sig00000db7,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ed7
    );
  blk00000001_blk00000ae8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dac,
      I1 => blk00000001_sig00000db8,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ed6
    );
  blk00000001_blk00000ae7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dad,
      I1 => blk00000001_sig00000db9,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ed5
    );
  blk00000001_blk00000ae6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dae,
      I1 => blk00000001_sig00000dba,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ed4
    );
  blk00000001_blk00000ae5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b9
    );
  blk00000001_blk00000ae4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001ba
    );
  blk00000001_blk00000ae3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001bf
    );
  blk00000001_blk00000ae2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ed0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001bb
    );
  blk00000001_blk00000ae1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd9,
      I1 => blk00000001_sig00000dca,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed3
    );
  blk00000001_blk00000ae0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dda,
      I1 => blk00000001_sig00000dcb,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed2
    );
  blk00000001_blk00000adf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000dd5,
      I1 => blk00000001_sig00000dcc,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed1
    );
  blk00000001_blk00000ade : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000ddb,
      I1 => blk00000001_sig00000dcd,
      I2 => blk00000001_sig00000dde,
      O => blk00000001_sig00000ed0
    );
  blk00000001_blk00000add : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ecf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c5
    );
  blk00000001_blk00000adc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ece,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c6
    );
  blk00000001_blk00000adb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ecd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c7
    );
  blk00000001_blk00000ada : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ecc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001c8
    );
  blk00000001_blk00000ad9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000da7,
      I1 => blk00000001_sig00000db7,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ecf
    );
  blk00000001_blk00000ad8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000da8,
      I1 => blk00000001_sig00000db8,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ece
    );
  blk00000001_blk00000ad7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000da9,
      I1 => blk00000001_sig00000db9,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ecd
    );
  blk00000001_blk00000ad6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000daa,
      I1 => blk00000001_sig00000dba,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000ecc
    );
  blk00000001_blk00000ad5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ecb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dda
    );
  blk00000001_blk00000ad4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eca,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000ddb
    );
  blk00000001_blk00000ad3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e98,
      I1 => blk00000001_sig00000e9b,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000ad3_O_UNCONNECTED
    );
  blk00000001_blk00000ad2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e97,
      I1 => blk00000001_sig00000e90,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ecb
    );
  blk00000001_blk00000ad1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e96,
      I1 => blk00000001_sig00000e99,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000ad1_O_UNCONNECTED
    );
  blk00000001_blk00000ad0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e95,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000eca
    );
  blk00000001_blk00000acf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd7
    );
  blk00000001_blk00000ace : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd8
    );
  blk00000001_blk00000acd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e89,
      I1 => blk00000001_sig00000e9b,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000acd_O_UNCONNECTED
    );
  blk00000001_blk00000acc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e8f,
      I1 => blk00000001_sig00000e8c,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec9
    );
  blk00000001_blk00000acb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e86,
      I1 => blk00000001_sig00000e99,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => NLW_blk00000001_blk00000acb_O_UNCONNECTED
    );
  blk00000001_blk00000aca : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e8e,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec8
    );
  blk00000001_blk00000ac9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd9
    );
  blk00000001_blk00000ac8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd4
    );
  blk00000001_blk00000ac7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd5
    );
  blk00000001_blk00000ac6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd6
    );
  blk00000001_blk00000ac5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e98,
      I1 => blk00000001_sig00000e9b,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec7
    );
  blk00000001_blk00000ac4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e88,
      I1 => blk00000001_sig00000e8d,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec6
    );
  blk00000001_blk00000ac3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e96,
      I1 => blk00000001_sig00000e99,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec5
    );
  blk00000001_blk00000ac2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e85,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec4
    );
  blk00000001_blk00000ac1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd0
    );
  blk00000001_blk00000ac0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd1
    );
  blk00000001_blk00000abf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd2
    );
  blk00000001_blk00000abe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ec0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dd3
    );
  blk00000001_blk00000abd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e89,
      I1 => blk00000001_sig00000e9b,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec3
    );
  blk00000001_blk00000abc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e8a,
      I1 => blk00000001_sig00000e8b,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec2
    );
  blk00000001_blk00000abb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e86,
      I1 => blk00000001_sig00000e99,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec1
    );
  blk00000001_blk00000aba : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000e87,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000ec0
    );
  blk00000001_blk00000ab9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ebf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e9f
    );
  blk00000001_blk00000ab8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ebe,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e9e
    );
  blk00000001_blk00000ab7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ebd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e9d
    );
  blk00000001_blk00000ab6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ebc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e9c
    );
  blk00000001_blk00000ab5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000eb2,
      I1 => blk00000001_sig00000ea8,
      I2 => blk00000001_sig00000eb2,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000ead,
      I5 => blk00000001_sig00000eae,
      O => blk00000001_sig00000ebf
    );
  blk00000001_blk00000ab4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000eb1,
      I1 => blk00000001_sig00000ea9,
      I2 => blk00000001_sig00000eb1,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000ead,
      I5 => blk00000001_sig00000eae,
      O => blk00000001_sig00000ebe
    );
  blk00000001_blk00000ab3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000ea8,
      I1 => blk00000001_sig00000eb0,
      I2 => blk00000001_sig00000eb0,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000ead,
      I5 => blk00000001_sig00000eae,
      O => blk00000001_sig00000ebd
    );
  blk00000001_blk00000ab2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000ea9,
      I1 => blk00000001_sig00000eaf,
      I2 => blk00000001_sig00000eaf,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000ead,
      I5 => blk00000001_sig00000eae,
      O => blk00000001_sig00000ebc
    );
  blk00000001_blk00000a9d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ebb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000ea7
    );
  blk00000001_blk00000a9c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eba,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000ea6
    );
  blk00000001_blk00000a9b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000ea9,
      Q => blk00000001_sig00000ebb
    );
  blk00000001_blk00000a9a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000ea8,
      Q => blk00000001_sig00000eba
    );
  blk00000001_blk00000a99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb9,
      Q => blk00000001_sig00000ea8
    );
  blk00000001_blk00000a98 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb8,
      Q => blk00000001_sig00000ea0
    );
  blk00000001_blk00000a97 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb7,
      Q => blk00000001_sig00000ea9
    );
  blk00000001_blk00000a96 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb6,
      Q => blk00000001_sig00000ea1
    );
  blk00000001_blk00000a95 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000eaa
    );
  blk00000001_blk00000a94 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dea,
      Q => blk00000001_sig00000eb5
    );
  blk00000001_blk00000a93 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000eac
    );
  blk00000001_blk00000a92 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000eb3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000eab
    );
  blk00000001_blk00000a91 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000e93,
      Q => blk00000001_sig00000eb4
    );
  blk00000001_blk00000a90 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000e94,
      Q => blk00000001_sig00000eb3
    );
  blk00000001_blk00000a8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000def,
      Q => blk00000001_sig00000eaf
    );
  blk00000001_blk00000a8e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000df0,
      Q => blk00000001_sig00000eb0
    );
  blk00000001_blk00000a8d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000df1,
      Q => blk00000001_sig00000eb1
    );
  blk00000001_blk00000a8c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000df2,
      Q => blk00000001_sig00000eb2
    );
  blk00000001_blk00000a8b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001b0,
      Q => blk00000001_sig00000ead
    );
  blk00000001_blk00000a8a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001b1,
      Q => blk00000001_sig00000eae
    );
  blk00000001_blk00000a89 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ea2,
      Q => blk00000001_sig00000e9b
    );
  blk00000001_blk00000a88 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ea3,
      Q => blk00000001_sig00000e9a
    );
  blk00000001_blk00000a87 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ea4,
      Q => blk00000001_sig00000e99
    );
  blk00000001_blk00000a86 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e9c,
      Q => blk00000001_sig00000e98
    );
  blk00000001_blk00000a85 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e9d,
      Q => blk00000001_sig00000e97
    );
  blk00000001_blk00000a84 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e9e,
      Q => blk00000001_sig00000e96
    );
  blk00000001_blk00000a83 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e9f,
      Q => blk00000001_sig00000e95
    );
  blk00000001_blk00000a82 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e84,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig0000009a
    );
  blk00000001_blk00000a81 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e83,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig00000099
    );
  blk00000001_blk00000a80 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e82,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig00000098
    );
  blk00000001_blk00000a7f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e81,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig00000097
    );
  blk00000001_blk00000a7e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e80,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig00000096
    );
  blk00000001_blk00000a7d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7f,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig00000095
    );
  blk00000001_blk00000a7c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df5,
      Q => blk00000001_sig00000e84
    );
  blk00000001_blk00000a7b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df6,
      Q => blk00000001_sig00000e83
    );
  blk00000001_blk00000a7a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df7,
      Q => blk00000001_sig00000e82
    );
  blk00000001_blk00000a79 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df8,
      Q => blk00000001_sig00000e81
    );
  blk00000001_blk00000a78 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df9,
      Q => blk00000001_sig00000e80
    );
  blk00000001_blk00000a77 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => blk00000001_sig000000c0,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dfa,
      Q => blk00000001_sig00000e7f
    );
  blk00000001_blk00000a76 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b5
    );
  blk00000001_blk00000a75 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b6
    );
  blk00000001_blk00000a74 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => blk00000001_sig000000c0,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001b7,
      Q => blk00000001_sig00000e7e
    );
  blk00000001_blk00000a73 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => blk00000001_sig000000c0,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001b8,
      Q => blk00000001_sig00000e7d
    );
  blk00000001_blk00000a60 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de1
    );
  blk00000001_blk00000a5f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de2
    );
  blk00000001_blk00000a5e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e7a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000a5e_Q_UNCONNECTED
    );
  blk00000001_blk00000a5d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001b0,
      Q => blk00000001_sig00000e7c
    );
  blk00000001_blk00000a5c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001b1,
      Q => blk00000001_sig00000e7b
    );
  blk00000001_blk00000a5b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001b2,
      Q => blk00000001_sig00000e7a
    );
  blk00000001_blk00000a5a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e79,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de3
    );
  blk00000001_blk00000a59 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e78,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de4
    );
  blk00000001_blk00000a58 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e77,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de5
    );
  blk00000001_blk00000a57 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e76,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000de6
    );
  blk00000001_blk00000a56 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000def,
      Q => blk00000001_sig00000e79
    );
  blk00000001_blk00000a55 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df0,
      Q => blk00000001_sig00000e78
    );
  blk00000001_blk00000a54 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df1,
      Q => blk00000001_sig00000e77
    );
  blk00000001_blk00000a53 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df2,
      Q => blk00000001_sig00000e76
    );
  blk00000001_blk00000a52 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e75,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000db7
    );
  blk00000001_blk00000a51 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e74,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000db8
    );
  blk00000001_blk00000a50 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e73,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000db9
    );
  blk00000001_blk00000a4f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e72,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000dba
    );
  blk00000001_blk00000a4e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dfd,
      Q => blk00000001_sig00000e75
    );
  blk00000001_blk00000a4d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dfe,
      Q => blk00000001_sig00000e74
    );
  blk00000001_blk00000a4c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dff,
      Q => blk00000001_sig00000e73
    );
  blk00000001_blk00000a4b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000e00,
      Q => blk00000001_sig00000e72
    );
  blk00000001_blk00000a4a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e71,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b7
    );
  blk00000001_blk00000a49 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e70,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b8
    );
  blk00000001_blk00000a48 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dce,
      Q => blk00000001_sig00000e71
    );
  blk00000001_blk00000a47 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dcf,
      Q => blk00000001_sig00000e70
    );
  blk00000001_blk00000a46 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e6f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b3
    );
  blk00000001_blk00000a45 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e6e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000001b4
    );
  blk00000001_blk00000a44 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df3,
      Q => blk00000001_sig00000e6f
    );
  blk00000001_blk00000a43 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000df4,
      Q => blk00000001_sig00000e6e
    );
  blk00000001_blk00000a14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0d,
      D => blk00000001_sig00000e6d,
      R => blk00000001_sig00000e12,
      Q => blk00000001_sig00000dea
    );
  blk00000001_blk00000a13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0d,
      D => blk00000001_sig00000e69,
      R => blk00000001_sig00000e12,
      Q => blk00000001_sig000001b2
    );
  blk00000001_blk00000a12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0d,
      D => blk00000001_sig00000e68,
      R => blk00000001_sig00000e12,
      Q => blk00000001_sig000001b1
    );
  blk00000001_blk00000a11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0d,
      D => blk00000001_sig00000e67,
      R => blk00000001_sig00000e12,
      Q => blk00000001_sig000001b0
    );
  blk00000001_blk000009fa : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000e61,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000e62,
      I3 => blk00000001_sig000000c0,
      I4 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e66
    );
  blk00000001_blk000009f9 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000e5e,
      I1 => blk00000001_sig000000c0,
      I2 => blk00000001_sig00000e5f,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000e60,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e65
    );
  blk00000001_blk000009f8 : MUXCY
    port map (
      CI => blk00000001_sig00000e63,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e66,
      O => blk00000001_sig00000e64
    );
  blk00000001_blk000009f7 : MUXCY
    port map (
      CI => blk00000001_sig000000c0,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e65,
      O => blk00000001_sig00000e63
    );
  blk00000001_blk000009f6 : XORCY
    port map (
      CI => blk00000001_sig00000e64,
      LI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e58
    );
  blk00000001_blk000009f5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e58,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e24
    );
  blk00000001_blk000009f4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e24,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig000001a8
    );
  blk00000001_blk000009f3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e57,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e62
    );
  blk00000001_blk000009f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e56,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e61
    );
  blk00000001_blk000009f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e55,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e60
    );
  blk00000001_blk000009f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e54,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e5f
    );
  blk00000001_blk000009ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0c,
      D => blk00000001_sig00000e53,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e5e
    );
  blk00000001_blk000009e1 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000df2,
      I1 => blk00000001_sig000000c0,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I5 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e52
    );
  blk00000001_blk000009e0 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000def,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000df0,
      I3 => blk00000001_sig000000c0,
      I4 => blk00000001_sig00000df1,
      I5 => blk00000001_sig000000c0,
      O => blk00000001_sig00000e51
    );
  blk00000001_blk000009df : MUXCY
    port map (
      CI => blk00000001_sig00000e4f,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e52,
      O => blk00000001_sig00000e50
    );
  blk00000001_blk000009de : MUXCY
    port map (
      CI => blk00000001_sig000000c0,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e51,
      O => blk00000001_sig00000e4f
    );
  blk00000001_blk000009dd : XORCY
    port map (
      CI => blk00000001_sig00000e50,
      LI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e4a
    );
  blk00000001_blk000009dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000deb,
      D => blk00000001_sig00000e4a,
      R => blk00000001_sig00000e0b,
      Q => blk00000001_sig00000e25
    );
  blk00000001_blk000009db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000deb,
      D => blk00000001_sig00000e49,
      R => blk00000001_sig00000e0b,
      Q => blk00000001_sig00000df2
    );
  blk00000001_blk000009da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000deb,
      D => blk00000001_sig00000e48,
      R => blk00000001_sig00000e0b,
      Q => blk00000001_sig00000df1
    );
  blk00000001_blk000009d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000deb,
      D => blk00000001_sig00000e47,
      R => blk00000001_sig00000e0b,
      Q => blk00000001_sig00000df0
    );
  blk00000001_blk000009d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000deb,
      D => blk00000001_sig00000e46,
      R => blk00000001_sig00000e0b,
      Q => blk00000001_sig00000def
    );
  blk00000001_blk000009c4 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000091,
      I1 => blk00000001_sig000000c0,
      I2 => blk00000001_sig00000090,
      I3 => blk00000001_sig000000c0,
      I4 => blk00000001_sig0000008f,
      I5 => blk00000001_sig000000c0,
      O => blk00000001_sig00000e45
    );
  blk00000001_blk000009c3 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig00000094,
      I1 => blk00000001_sig000000c0,
      I2 => blk00000001_sig00000093,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig00000092,
      I5 => blk00000001_sig000000c0,
      O => blk00000001_sig00000e44
    );
  blk00000001_blk000009c2 : MUXCY
    port map (
      CI => blk00000001_sig00000e42,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e45,
      O => blk00000001_sig00000e43
    );
  blk00000001_blk000009c1 : MUXCY
    port map (
      CI => blk00000001_sig000000c0,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig00000e44,
      O => blk00000001_sig00000e42
    );
  blk00000001_blk000009c0 : XORCY
    port map (
      CI => blk00000001_sig00000e43,
      LI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      O => blk00000001_sig00000e3b
    );
  blk00000001_blk000009bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e3b,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e27
    );
  blk00000001_blk000009be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e27,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e26
    );
  blk00000001_blk000009bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e3a,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig0000008f
    );
  blk00000001_blk000009bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e39,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000090
    );
  blk00000001_blk000009bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e38,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000091
    );
  blk00000001_blk000009ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e37,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000092
    );
  blk00000001_blk000009b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e36,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000093
    );
  blk00000001_blk000009b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig00000e0e,
      D => blk00000001_sig00000e35,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000094
    );
  blk00000001_blk000009b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e09,
      Q => blk00000001_sig000001a4
    );
  blk00000001_blk000009b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e03,
      Q => blk00000001_sig00000e17
    );
  blk00000001_blk000009b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e04,
      Q => blk00000001_sig00000e18
    );
  blk00000001_blk000009b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e06,
      Q => blk00000001_sig00000e19
    );
  blk00000001_blk000009b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e05,
      Q => blk00000001_sig00000e1a
    );
  blk00000001_blk000009b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e0a,
      Q => blk00000001_sig00000de9
    );
  blk00000001_blk000009b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e08,
      Q => blk00000001_sig00000e14
    );
  blk00000001_blk000009b0 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e07,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e0f
    );
  blk00000001_blk000009af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000090,
      Q => blk00000001_sig00000dfd
    );
  blk00000001_blk000009ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000008f,
      Q => blk00000001_sig00000dfe
    );
  blk00000001_blk000009ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000092,
      Q => blk00000001_sig00000dff
    );
  blk00000001_blk000009ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000091,
      Q => blk00000001_sig00000e00
    );
  blk00000001_blk000009ab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000bb,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e11
    );
  blk00000001_blk000009aa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e16,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000e10
    );
  blk00000001_blk000009a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000094,
      Q => blk00000001_sig00000dfb
    );
  blk00000001_blk000009a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000093,
      Q => blk00000001_sig00000dfc
    );
  blk00000001_blk000009a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e23,
      Q => blk00000001_sig00000e1d
    );
  blk00000001_blk000009a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e02,
      Q => blk00000001_sig00000e1b
    );
  blk00000001_blk000009a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e01,
      Q => blk00000001_sig00000e1c
    );
  blk00000001_blk000009a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e1b,
      Q => blk00000001_sig00000df3
    );
  blk00000001_blk000009a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000e1c,
      Q => blk00000001_sig00000df4
    );
  blk00000001_blk000009a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e34
    );
  blk00000001_blk000009a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e33
    );
  blk00000001_blk000009a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e32
    );
  blk00000001_blk0000099f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e31
    );
  blk00000001_blk0000099e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e30
    );
  blk00000001_blk0000099d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2f
    );
  blk00000001_blk0000099c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2e
    );
  blk00000001_blk0000099b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2d
    );
  blk00000001_blk0000099a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2c
    );
  blk00000001_blk00000999 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2b
    );
  blk00000001_blk00000998 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e2a
    );
  blk00000001_blk00000997 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000e29
    );
  blk00000001_blk00000996 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000c0,
      Q => blk00000001_sig00000e28
    );
  blk00000001_blk00000995 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da5,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig000001a7
    );
  blk00000001_blk00000994 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da1,
      Q => blk00000001_sig000001d5
    );
  blk00000001_blk00000993 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da2,
      Q => blk00000001_sig000001d6
    );
  blk00000001_blk00000992 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da3,
      Q => blk00000001_sig000001d7
    );
  blk00000001_blk00000991 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da4,
      Q => blk00000001_sig000001d8
    );
  blk00000001_blk00000990 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000dee,
      Q => blk00000001_sig00000ddd
    );
  blk00000001_blk000008e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d1
    );
  blk00000001_blk000008e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d2
    );
  blk00000001_blk000008e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d3
    );
  blk00000001_blk000008e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d4
    );
  blk00000001_blk000008e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d5
    );
  blk00000001_blk000008e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d6
    );
  blk00000001_blk000008df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d9a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d7
    );
  blk00000001_blk000008de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d99,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d8
    );
  blk00000001_blk000008dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d98,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d9
    );
  blk00000001_blk000008dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d97,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002da
    );
  blk00000001_blk000008db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d96,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002db
    );
  blk00000001_blk000008da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d95,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002dc
    );
  blk00000001_blk000008d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d94,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002dd
    );
  blk00000001_blk000008d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d93,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002de
    );
  blk00000001_blk000008d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d92,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002df
    );
  blk00000001_blk000008d6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d91,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e0
    );
  blk00000001_blk000008d5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000327,
      I1 => blk00000001_sig0000041e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000da0
    );
  blk00000001_blk000008d4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000328,
      I1 => blk00000001_sig0000041f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9f
    );
  blk00000001_blk000008d3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000329,
      I1 => blk00000001_sig00000420,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9e
    );
  blk00000001_blk000008d2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032a,
      I1 => blk00000001_sig00000421,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9d
    );
  blk00000001_blk000008d1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032b,
      I1 => blk00000001_sig00000422,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9c
    );
  blk00000001_blk000008d0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032c,
      I1 => blk00000001_sig00000423,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9b
    );
  blk00000001_blk000008cf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032d,
      I1 => blk00000001_sig00000424,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d9a
    );
  blk00000001_blk000008ce : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032e,
      I1 => blk00000001_sig00000425,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d99
    );
  blk00000001_blk000008cd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000032f,
      I1 => blk00000001_sig00000426,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d98
    );
  blk00000001_blk000008cc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000330,
      I1 => blk00000001_sig00000427,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d97
    );
  blk00000001_blk000008cb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000331,
      I1 => blk00000001_sig00000428,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d96
    );
  blk00000001_blk000008ca : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000332,
      I1 => blk00000001_sig00000429,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d95
    );
  blk00000001_blk000008c9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000333,
      I1 => blk00000001_sig0000042a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d94
    );
  blk00000001_blk000008c8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000334,
      I1 => blk00000001_sig0000042b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d93
    );
  blk00000001_blk000008c7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000335,
      I1 => blk00000001_sig0000042c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d92
    );
  blk00000001_blk000008c6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000336,
      I1 => blk00000001_sig0000042d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d91
    );
  blk00000001_blk000008c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d90,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c1
    );
  blk00000001_blk000008c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c2
    );
  blk00000001_blk000008c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c3
    );
  blk00000001_blk000008c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c4
    );
  blk00000001_blk000008c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c5
    );
  blk00000001_blk000008c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c6
    );
  blk00000001_blk000008bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d8a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c7
    );
  blk00000001_blk000008be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d89,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c8
    );
  blk00000001_blk000008bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d88,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c9
    );
  blk00000001_blk000008bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d87,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ca
    );
  blk00000001_blk000008bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d86,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002cb
    );
  blk00000001_blk000008ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d85,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002cc
    );
  blk00000001_blk000008b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d84,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002cd
    );
  blk00000001_blk000008b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d83,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ce
    );
  blk00000001_blk000008b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d82,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002cf
    );
  blk00000001_blk000008b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d81,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002d0
    );
  blk00000001_blk000008b5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002e7,
      I1 => blk00000001_sig0000040e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d90
    );
  blk00000001_blk000008b4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002e8,
      I1 => blk00000001_sig0000040f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8f
    );
  blk00000001_blk000008b3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002e9,
      I1 => blk00000001_sig00000410,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8e
    );
  blk00000001_blk000008b2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ea,
      I1 => blk00000001_sig00000411,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8d
    );
  blk00000001_blk000008b1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002eb,
      I1 => blk00000001_sig00000412,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8c
    );
  blk00000001_blk000008b0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ec,
      I1 => blk00000001_sig00000413,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8b
    );
  blk00000001_blk000008af : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ed,
      I1 => blk00000001_sig00000414,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d8a
    );
  blk00000001_blk000008ae : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ee,
      I1 => blk00000001_sig00000415,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d89
    );
  blk00000001_blk000008ad : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ef,
      I1 => blk00000001_sig00000416,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d88
    );
  blk00000001_blk000008ac : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f0,
      I1 => blk00000001_sig00000417,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d87
    );
  blk00000001_blk000008ab : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f1,
      I1 => blk00000001_sig00000418,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d86
    );
  blk00000001_blk000008aa : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f2,
      I1 => blk00000001_sig00000419,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d85
    );
  blk00000001_blk000008a9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f3,
      I1 => blk00000001_sig0000041a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d84
    );
  blk00000001_blk000008a8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f4,
      I1 => blk00000001_sig0000041b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d83
    );
  blk00000001_blk000008a7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f5,
      I1 => blk00000001_sig0000041c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d82
    );
  blk00000001_blk000008a6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f6,
      I1 => blk00000001_sig0000041d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d81
    );
  blk00000001_blk000008a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d80,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b1
    );
  blk00000001_blk000008a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b2
    );
  blk00000001_blk000008a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b3
    );
  blk00000001_blk000008a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b4
    );
  blk00000001_blk000008a1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b5
    );
  blk00000001_blk000008a0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b6
    );
  blk00000001_blk0000089f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d7a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b7
    );
  blk00000001_blk0000089e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d79,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b8
    );
  blk00000001_blk0000089d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d78,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b9
    );
  blk00000001_blk0000089c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d77,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ba
    );
  blk00000001_blk0000089b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d76,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002bb
    );
  blk00000001_blk0000089a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d75,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002bc
    );
  blk00000001_blk00000899 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d74,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002bd
    );
  blk00000001_blk00000898 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d73,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002be
    );
  blk00000001_blk00000897 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d72,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002bf
    );
  blk00000001_blk00000896 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d71,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002c0
    );
  blk00000001_blk00000895 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000337,
      I1 => blk00000001_sig0000041e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d80
    );
  blk00000001_blk00000894 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000338,
      I1 => blk00000001_sig0000041f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7f
    );
  blk00000001_blk00000893 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000339,
      I1 => blk00000001_sig00000420,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7e
    );
  blk00000001_blk00000892 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033a,
      I1 => blk00000001_sig00000421,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7d
    );
  blk00000001_blk00000891 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033b,
      I1 => blk00000001_sig00000422,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7c
    );
  blk00000001_blk00000890 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033c,
      I1 => blk00000001_sig00000423,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7b
    );
  blk00000001_blk0000088f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033d,
      I1 => blk00000001_sig00000424,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d7a
    );
  blk00000001_blk0000088e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033e,
      I1 => blk00000001_sig00000425,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d79
    );
  blk00000001_blk0000088d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000033f,
      I1 => blk00000001_sig00000426,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d78
    );
  blk00000001_blk0000088c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000340,
      I1 => blk00000001_sig00000427,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d77
    );
  blk00000001_blk0000088b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000341,
      I1 => blk00000001_sig00000428,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d76
    );
  blk00000001_blk0000088a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000342,
      I1 => blk00000001_sig00000429,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d75
    );
  blk00000001_blk00000889 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000343,
      I1 => blk00000001_sig0000042a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d74
    );
  blk00000001_blk00000888 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000344,
      I1 => blk00000001_sig0000042b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d73
    );
  blk00000001_blk00000887 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000345,
      I1 => blk00000001_sig0000042c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d72
    );
  blk00000001_blk00000886 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000346,
      I1 => blk00000001_sig0000042d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d71
    );
  blk00000001_blk00000885 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d70,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a1
    );
  blk00000001_blk00000884 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a2
    );
  blk00000001_blk00000883 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a3
    );
  blk00000001_blk00000882 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a4
    );
  blk00000001_blk00000881 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a5
    );
  blk00000001_blk00000880 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a6
    );
  blk00000001_blk0000087f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d6a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a7
    );
  blk00000001_blk0000087e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d69,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a8
    );
  blk00000001_blk0000087d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d68,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a9
    );
  blk00000001_blk0000087c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d67,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002aa
    );
  blk00000001_blk0000087b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d66,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ab
    );
  blk00000001_blk0000087a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d65,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ac
    );
  blk00000001_blk00000879 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d64,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ad
    );
  blk00000001_blk00000878 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d63,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ae
    );
  blk00000001_blk00000877 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d62,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002af
    );
  blk00000001_blk00000876 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d61,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002b0
    );
  blk00000001_blk00000875 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f7,
      I1 => blk00000001_sig0000040e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d70
    );
  blk00000001_blk00000874 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f8,
      I1 => blk00000001_sig0000040f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6f
    );
  blk00000001_blk00000873 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002f9,
      I1 => blk00000001_sig00000410,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6e
    );
  blk00000001_blk00000872 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002fa,
      I1 => blk00000001_sig00000411,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6d
    );
  blk00000001_blk00000871 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002fb,
      I1 => blk00000001_sig00000412,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6c
    );
  blk00000001_blk00000870 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002fc,
      I1 => blk00000001_sig00000413,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6b
    );
  blk00000001_blk0000086f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002fd,
      I1 => blk00000001_sig00000414,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d6a
    );
  blk00000001_blk0000086e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002fe,
      I1 => blk00000001_sig00000415,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d69
    );
  blk00000001_blk0000086d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig000002ff,
      I1 => blk00000001_sig00000416,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d68
    );
  blk00000001_blk0000086c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000300,
      I1 => blk00000001_sig00000417,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d67
    );
  blk00000001_blk0000086b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000301,
      I1 => blk00000001_sig00000418,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d66
    );
  blk00000001_blk0000086a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000302,
      I1 => blk00000001_sig00000419,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d65
    );
  blk00000001_blk00000869 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000303,
      I1 => blk00000001_sig0000041a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d64
    );
  blk00000001_blk00000868 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000304,
      I1 => blk00000001_sig0000041b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d63
    );
  blk00000001_blk00000867 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000305,
      I1 => blk00000001_sig0000041c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d62
    );
  blk00000001_blk00000866 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000306,
      I1 => blk00000001_sig0000041d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d61
    );
  blk00000001_blk00000865 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d60,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000291
    );
  blk00000001_blk00000864 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000292
    );
  blk00000001_blk00000863 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000293
    );
  blk00000001_blk00000862 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000294
    );
  blk00000001_blk00000861 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000295
    );
  blk00000001_blk00000860 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000296
    );
  blk00000001_blk0000085f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d5a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000297
    );
  blk00000001_blk0000085e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d59,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000298
    );
  blk00000001_blk0000085d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d58,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000299
    );
  blk00000001_blk0000085c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d57,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029a
    );
  blk00000001_blk0000085b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d56,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029b
    );
  blk00000001_blk0000085a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d55,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029c
    );
  blk00000001_blk00000859 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d54,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029d
    );
  blk00000001_blk00000858 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d53,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029e
    );
  blk00000001_blk00000857 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d52,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000029f
    );
  blk00000001_blk00000856 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d51,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002a0
    );
  blk00000001_blk00000855 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000347,
      I1 => blk00000001_sig0000041e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d60
    );
  blk00000001_blk00000854 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000348,
      I1 => blk00000001_sig0000041f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5f
    );
  blk00000001_blk00000853 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000349,
      I1 => blk00000001_sig00000420,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5e
    );
  blk00000001_blk00000852 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034a,
      I1 => blk00000001_sig00000421,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5d
    );
  blk00000001_blk00000851 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034b,
      I1 => blk00000001_sig00000422,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5c
    );
  blk00000001_blk00000850 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034c,
      I1 => blk00000001_sig00000423,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5b
    );
  blk00000001_blk0000084f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034d,
      I1 => blk00000001_sig00000424,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d5a
    );
  blk00000001_blk0000084e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034e,
      I1 => blk00000001_sig00000425,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d59
    );
  blk00000001_blk0000084d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000034f,
      I1 => blk00000001_sig00000426,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d58
    );
  blk00000001_blk0000084c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000350,
      I1 => blk00000001_sig00000427,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d57
    );
  blk00000001_blk0000084b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000351,
      I1 => blk00000001_sig00000428,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d56
    );
  blk00000001_blk0000084a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000352,
      I1 => blk00000001_sig00000429,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d55
    );
  blk00000001_blk00000849 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000353,
      I1 => blk00000001_sig0000042a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d54
    );
  blk00000001_blk00000848 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000354,
      I1 => blk00000001_sig0000042b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d53
    );
  blk00000001_blk00000847 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000355,
      I1 => blk00000001_sig0000042c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d52
    );
  blk00000001_blk00000846 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000356,
      I1 => blk00000001_sig0000042d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d51
    );
  blk00000001_blk00000845 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d50,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000281
    );
  blk00000001_blk00000844 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000282
    );
  blk00000001_blk00000843 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000283
    );
  blk00000001_blk00000842 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000284
    );
  blk00000001_blk00000841 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000285
    );
  blk00000001_blk00000840 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000286
    );
  blk00000001_blk0000083f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d4a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000287
    );
  blk00000001_blk0000083e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d49,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000288
    );
  blk00000001_blk0000083d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d48,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000289
    );
  blk00000001_blk0000083c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d47,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028a
    );
  blk00000001_blk0000083b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d46,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028b
    );
  blk00000001_blk0000083a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d45,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028c
    );
  blk00000001_blk00000839 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d44,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028d
    );
  blk00000001_blk00000838 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d43,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028e
    );
  blk00000001_blk00000837 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d42,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000028f
    );
  blk00000001_blk00000836 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d41,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000290
    );
  blk00000001_blk00000835 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000307,
      I1 => blk00000001_sig0000040e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d50
    );
  blk00000001_blk00000834 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000308,
      I1 => blk00000001_sig0000040f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4f
    );
  blk00000001_blk00000833 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000309,
      I1 => blk00000001_sig00000410,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4e
    );
  blk00000001_blk00000832 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030a,
      I1 => blk00000001_sig00000411,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4d
    );
  blk00000001_blk00000831 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030b,
      I1 => blk00000001_sig00000412,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4c
    );
  blk00000001_blk00000830 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030c,
      I1 => blk00000001_sig00000413,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4b
    );
  blk00000001_blk0000082f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030d,
      I1 => blk00000001_sig00000414,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d4a
    );
  blk00000001_blk0000082e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030e,
      I1 => blk00000001_sig00000415,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d49
    );
  blk00000001_blk0000082d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000030f,
      I1 => blk00000001_sig00000416,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d48
    );
  blk00000001_blk0000082c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000310,
      I1 => blk00000001_sig00000417,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d47
    );
  blk00000001_blk0000082b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000311,
      I1 => blk00000001_sig00000418,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d46
    );
  blk00000001_blk0000082a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000312,
      I1 => blk00000001_sig00000419,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d45
    );
  blk00000001_blk00000829 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000313,
      I1 => blk00000001_sig0000041a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d44
    );
  blk00000001_blk00000828 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000314,
      I1 => blk00000001_sig0000041b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d43
    );
  blk00000001_blk00000827 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000315,
      I1 => blk00000001_sig0000041c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d42
    );
  blk00000001_blk00000826 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000316,
      I1 => blk00000001_sig0000041d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d41
    );
  blk00000001_blk00000825 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d40,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000271
    );
  blk00000001_blk00000824 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000272
    );
  blk00000001_blk00000823 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000273
    );
  blk00000001_blk00000822 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000274
    );
  blk00000001_blk00000821 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000275
    );
  blk00000001_blk00000820 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000276
    );
  blk00000001_blk0000081f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d3a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000277
    );
  blk00000001_blk0000081e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d39,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000278
    );
  blk00000001_blk0000081d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d38,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000279
    );
  blk00000001_blk0000081c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d37,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027a
    );
  blk00000001_blk0000081b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d36,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027b
    );
  blk00000001_blk0000081a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d35,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027c
    );
  blk00000001_blk00000819 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d34,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027d
    );
  blk00000001_blk00000818 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d33,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027e
    );
  blk00000001_blk00000817 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d32,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000027f
    );
  blk00000001_blk00000816 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d31,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000280
    );
  blk00000001_blk00000815 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000357,
      I1 => blk00000001_sig0000041e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d40
    );
  blk00000001_blk00000814 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000358,
      I1 => blk00000001_sig0000041f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3f
    );
  blk00000001_blk00000813 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000359,
      I1 => blk00000001_sig00000420,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3e
    );
  blk00000001_blk00000812 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035a,
      I1 => blk00000001_sig00000421,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3d
    );
  blk00000001_blk00000811 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035b,
      I1 => blk00000001_sig00000422,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3c
    );
  blk00000001_blk00000810 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035c,
      I1 => blk00000001_sig00000423,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3b
    );
  blk00000001_blk0000080f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035d,
      I1 => blk00000001_sig00000424,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d3a
    );
  blk00000001_blk0000080e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035e,
      I1 => blk00000001_sig00000425,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d39
    );
  blk00000001_blk0000080d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000035f,
      I1 => blk00000001_sig00000426,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d38
    );
  blk00000001_blk0000080c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000360,
      I1 => blk00000001_sig00000427,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d37
    );
  blk00000001_blk0000080b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000361,
      I1 => blk00000001_sig00000428,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d36
    );
  blk00000001_blk0000080a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000362,
      I1 => blk00000001_sig00000429,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d35
    );
  blk00000001_blk00000809 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000363,
      I1 => blk00000001_sig0000042a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d34
    );
  blk00000001_blk00000808 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000364,
      I1 => blk00000001_sig0000042b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d33
    );
  blk00000001_blk00000807 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000365,
      I1 => blk00000001_sig0000042c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d32
    );
  blk00000001_blk00000806 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000366,
      I1 => blk00000001_sig0000042d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d31
    );
  blk00000001_blk00000805 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d30,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000261
    );
  blk00000001_blk00000804 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000262
    );
  blk00000001_blk00000803 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000263
    );
  blk00000001_blk00000802 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000264
    );
  blk00000001_blk00000801 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000265
    );
  blk00000001_blk00000800 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000266
    );
  blk00000001_blk000007ff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d2a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000267
    );
  blk00000001_blk000007fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d29,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000268
    );
  blk00000001_blk000007fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d28,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000269
    );
  blk00000001_blk000007fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d27,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026a
    );
  blk00000001_blk000007fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d26,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026b
    );
  blk00000001_blk000007fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d25,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026c
    );
  blk00000001_blk000007f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d24,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026d
    );
  blk00000001_blk000007f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d23,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026e
    );
  blk00000001_blk000007f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d22,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000026f
    );
  blk00000001_blk000007f6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d21,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000270
    );
  blk00000001_blk000007f5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000317,
      I1 => blk00000001_sig0000040e,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d30
    );
  blk00000001_blk000007f4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000318,
      I1 => blk00000001_sig0000040f,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2f
    );
  blk00000001_blk000007f3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000319,
      I1 => blk00000001_sig00000410,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2e
    );
  blk00000001_blk000007f2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031a,
      I1 => blk00000001_sig00000411,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2d
    );
  blk00000001_blk000007f1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031b,
      I1 => blk00000001_sig00000412,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2c
    );
  blk00000001_blk000007f0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031c,
      I1 => blk00000001_sig00000413,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2b
    );
  blk00000001_blk000007ef : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031d,
      I1 => blk00000001_sig00000414,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d2a
    );
  blk00000001_blk000007ee : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031e,
      I1 => blk00000001_sig00000415,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d29
    );
  blk00000001_blk000007ed : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig0000031f,
      I1 => blk00000001_sig00000416,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d28
    );
  blk00000001_blk000007ec : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000320,
      I1 => blk00000001_sig00000417,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d27
    );
  blk00000001_blk000007eb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000321,
      I1 => blk00000001_sig00000418,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d26
    );
  blk00000001_blk000007ea : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000322,
      I1 => blk00000001_sig00000419,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d25
    );
  blk00000001_blk000007e9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000323,
      I1 => blk00000001_sig0000041a,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d24
    );
  blk00000001_blk000007e8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000324,
      I1 => blk00000001_sig0000041b,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d23
    );
  blk00000001_blk000007e7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000325,
      I1 => blk00000001_sig0000041c,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d22
    );
  blk00000001_blk000007e6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_sig00000326,
      I1 => blk00000001_sig0000041d,
      I2 => blk00000001_sig000001af,
      O => blk00000001_sig00000d21
    );
  blk00000001_blk000007df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d1c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e6
    );
  blk00000001_blk000007de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d1b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e5
    );
  blk00000001_blk000007dd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001db,
      I1 => blk00000001_sig000001dd,
      I2 => blk00000001_sig000001df,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig000001b0,
      I5 => blk00000001_sig000001b1,
      O => blk00000001_sig00000d20
    );
  blk00000001_blk000007dc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001da,
      I1 => blk00000001_sig000001dc,
      I2 => blk00000001_sig000001de,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig000001b0,
      I5 => blk00000001_sig000001b1,
      O => blk00000001_sig00000d1f
    );
  blk00000001_blk000007db : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig000001b0,
      I5 => blk00000001_sig000001b1,
      O => blk00000001_sig00000d1e
    );
  blk00000001_blk000007da : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I4 => blk00000001_sig000001b0,
      I5 => blk00000001_sig000001b1,
      O => blk00000001_sig00000d1d
    );
  blk00000001_blk000007d9 : MUXF7
    port map (
      I0 => blk00000001_sig00000d20,
      I1 => blk00000001_sig00000d1e,
      S => blk00000001_sig000001b2,
      O => blk00000001_sig00000d1c
    );
  blk00000001_blk000007d8 : MUXF7
    port map (
      I0 => blk00000001_sig00000d1f,
      I1 => blk00000001_sig00000d1d,
      S => blk00000001_sig000001b2,
      O => blk00000001_sig00000d1b
    );
  blk00000001_blk000007d7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d8,
      I1 => blk00000001_sig000003b8,
      I2 => blk00000001_sig00000398,
      I3 => blk00000001_sig00000378,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d1a
    );
  blk00000001_blk000007d6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d9,
      I1 => blk00000001_sig000003b9,
      I2 => blk00000001_sig00000399,
      I3 => blk00000001_sig00000379,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d19
    );
  blk00000001_blk000007d5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003da,
      I1 => blk00000001_sig000003ba,
      I2 => blk00000001_sig0000039a,
      I3 => blk00000001_sig0000037a,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d18
    );
  blk00000001_blk000007d4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003db,
      I1 => blk00000001_sig000003bb,
      I2 => blk00000001_sig0000039b,
      I3 => blk00000001_sig0000037b,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d17
    );
  blk00000001_blk000007d3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dc,
      I1 => blk00000001_sig000003bc,
      I2 => blk00000001_sig0000039c,
      I3 => blk00000001_sig0000037c,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d16
    );
  blk00000001_blk000007d2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dd,
      I1 => blk00000001_sig000003bd,
      I2 => blk00000001_sig0000039d,
      I3 => blk00000001_sig0000037d,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d15
    );
  blk00000001_blk000007d1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003de,
      I1 => blk00000001_sig000003be,
      I2 => blk00000001_sig0000039e,
      I3 => blk00000001_sig0000037e,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d14
    );
  blk00000001_blk000007d0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003df,
      I1 => blk00000001_sig000003bf,
      I2 => blk00000001_sig0000039f,
      I3 => blk00000001_sig0000037f,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d13
    );
  blk00000001_blk000007cf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e0,
      I1 => blk00000001_sig000003c0,
      I2 => blk00000001_sig000003a0,
      I3 => blk00000001_sig00000380,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d12
    );
  blk00000001_blk000007ce : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e1,
      I1 => blk00000001_sig000003c1,
      I2 => blk00000001_sig000003a1,
      I3 => blk00000001_sig00000381,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d11
    );
  blk00000001_blk000007cd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e2,
      I1 => blk00000001_sig000003c2,
      I2 => blk00000001_sig000003a2,
      I3 => blk00000001_sig00000382,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d10
    );
  blk00000001_blk000007cc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e3,
      I1 => blk00000001_sig000003c3,
      I2 => blk00000001_sig000003a3,
      I3 => blk00000001_sig00000383,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d0f
    );
  blk00000001_blk000007cb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e4,
      I1 => blk00000001_sig000003c4,
      I2 => blk00000001_sig000003a4,
      I3 => blk00000001_sig00000384,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d0e
    );
  blk00000001_blk000007ca : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e5,
      I1 => blk00000001_sig000003c5,
      I2 => blk00000001_sig000003a5,
      I3 => blk00000001_sig00000385,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d0d
    );
  blk00000001_blk000007c9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e6,
      I1 => blk00000001_sig000003c6,
      I2 => blk00000001_sig000003a6,
      I3 => blk00000001_sig00000386,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d0c
    );
  blk00000001_blk000007c8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e7,
      I1 => blk00000001_sig000003c7,
      I2 => blk00000001_sig000003a7,
      I3 => blk00000001_sig00000387,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000d0b
    );
  blk00000001_blk000007c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d1a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000327
    );
  blk00000001_blk000007c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d19,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000328
    );
  blk00000001_blk000007c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d18,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000329
    );
  blk00000001_blk000007c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d17,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032a
    );
  blk00000001_blk000007c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d16,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032b
    );
  blk00000001_blk000007c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d15,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032c
    );
  blk00000001_blk000007c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d14,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032d
    );
  blk00000001_blk000007c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d13,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032e
    );
  blk00000001_blk000007bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d12,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000032f
    );
  blk00000001_blk000007be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d11,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000330
    );
  blk00000001_blk000007bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d10,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000331
    );
  blk00000001_blk000007bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000332
    );
  blk00000001_blk000007bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000333
    );
  blk00000001_blk000007ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000334
    );
  blk00000001_blk000007b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000335
    );
  blk00000001_blk000007b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000336
    );
  blk00000001_blk000007b7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d8,
      I1 => blk00000001_sig000003b8,
      I2 => blk00000001_sig00000398,
      I3 => blk00000001_sig00000378,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d0a
    );
  blk00000001_blk000007b6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d9,
      I1 => blk00000001_sig000003b9,
      I2 => blk00000001_sig00000399,
      I3 => blk00000001_sig00000379,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d09
    );
  blk00000001_blk000007b5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003da,
      I1 => blk00000001_sig000003ba,
      I2 => blk00000001_sig0000039a,
      I3 => blk00000001_sig0000037a,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d08
    );
  blk00000001_blk000007b4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003db,
      I1 => blk00000001_sig000003bb,
      I2 => blk00000001_sig0000039b,
      I3 => blk00000001_sig0000037b,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d07
    );
  blk00000001_blk000007b3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dc,
      I1 => blk00000001_sig000003bc,
      I2 => blk00000001_sig0000039c,
      I3 => blk00000001_sig0000037c,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d06
    );
  blk00000001_blk000007b2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dd,
      I1 => blk00000001_sig000003bd,
      I2 => blk00000001_sig0000039d,
      I3 => blk00000001_sig0000037d,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d05
    );
  blk00000001_blk000007b1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003de,
      I1 => blk00000001_sig000003be,
      I2 => blk00000001_sig0000039e,
      I3 => blk00000001_sig0000037e,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d04
    );
  blk00000001_blk000007b0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003df,
      I1 => blk00000001_sig000003bf,
      I2 => blk00000001_sig0000039f,
      I3 => blk00000001_sig0000037f,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d03
    );
  blk00000001_blk000007af : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e0,
      I1 => blk00000001_sig000003c0,
      I2 => blk00000001_sig000003a0,
      I3 => blk00000001_sig00000380,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d02
    );
  blk00000001_blk000007ae : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e1,
      I1 => blk00000001_sig000003c1,
      I2 => blk00000001_sig000003a1,
      I3 => blk00000001_sig00000381,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d01
    );
  blk00000001_blk000007ad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e2,
      I1 => blk00000001_sig000003c2,
      I2 => blk00000001_sig000003a2,
      I3 => blk00000001_sig00000382,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000d00
    );
  blk00000001_blk000007ac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e3,
      I1 => blk00000001_sig000003c3,
      I2 => blk00000001_sig000003a3,
      I3 => blk00000001_sig00000383,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cff
    );
  blk00000001_blk000007ab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e4,
      I1 => blk00000001_sig000003c4,
      I2 => blk00000001_sig000003a4,
      I3 => blk00000001_sig00000384,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cfe
    );
  blk00000001_blk000007aa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e5,
      I1 => blk00000001_sig000003c5,
      I2 => blk00000001_sig000003a5,
      I3 => blk00000001_sig00000385,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cfd
    );
  blk00000001_blk000007a9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e6,
      I1 => blk00000001_sig000003c6,
      I2 => blk00000001_sig000003a6,
      I3 => blk00000001_sig00000386,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cfc
    );
  blk00000001_blk000007a8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e7,
      I1 => blk00000001_sig000003c7,
      I2 => blk00000001_sig000003a7,
      I3 => blk00000001_sig00000387,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cfb
    );
  blk00000001_blk000007a7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d0a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000337
    );
  blk00000001_blk000007a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d09,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000338
    );
  blk00000001_blk000007a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d08,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000339
    );
  blk00000001_blk000007a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d07,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033a
    );
  blk00000001_blk000007a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d06,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033b
    );
  blk00000001_blk000007a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d05,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033c
    );
  blk00000001_blk000007a1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d04,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033d
    );
  blk00000001_blk000007a0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d03,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033e
    );
  blk00000001_blk0000079f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d02,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000033f
    );
  blk00000001_blk0000079e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d01,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000340
    );
  blk00000001_blk0000079d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000d00,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000341
    );
  blk00000001_blk0000079c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cff,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000342
    );
  blk00000001_blk0000079b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cfe,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000343
    );
  blk00000001_blk0000079a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cfd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000344
    );
  blk00000001_blk00000799 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cfc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000345
    );
  blk00000001_blk00000798 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cfb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000346
    );
  blk00000001_blk00000797 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d8,
      I1 => blk00000001_sig000003b8,
      I2 => blk00000001_sig00000398,
      I3 => blk00000001_sig00000378,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cfa
    );
  blk00000001_blk00000796 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d9,
      I1 => blk00000001_sig000003b9,
      I2 => blk00000001_sig00000399,
      I3 => blk00000001_sig00000379,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf9
    );
  blk00000001_blk00000795 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003da,
      I1 => blk00000001_sig000003ba,
      I2 => blk00000001_sig0000039a,
      I3 => blk00000001_sig0000037a,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf8
    );
  blk00000001_blk00000794 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003db,
      I1 => blk00000001_sig000003bb,
      I2 => blk00000001_sig0000039b,
      I3 => blk00000001_sig0000037b,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf7
    );
  blk00000001_blk00000793 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dc,
      I1 => blk00000001_sig000003bc,
      I2 => blk00000001_sig0000039c,
      I3 => blk00000001_sig0000037c,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf6
    );
  blk00000001_blk00000792 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dd,
      I1 => blk00000001_sig000003bd,
      I2 => blk00000001_sig0000039d,
      I3 => blk00000001_sig0000037d,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf5
    );
  blk00000001_blk00000791 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003de,
      I1 => blk00000001_sig000003be,
      I2 => blk00000001_sig0000039e,
      I3 => blk00000001_sig0000037e,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf4
    );
  blk00000001_blk00000790 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003df,
      I1 => blk00000001_sig000003bf,
      I2 => blk00000001_sig0000039f,
      I3 => blk00000001_sig0000037f,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf3
    );
  blk00000001_blk0000078f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e0,
      I1 => blk00000001_sig000003c0,
      I2 => blk00000001_sig000003a0,
      I3 => blk00000001_sig00000380,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf2
    );
  blk00000001_blk0000078e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e1,
      I1 => blk00000001_sig000003c1,
      I2 => blk00000001_sig000003a1,
      I3 => blk00000001_sig00000381,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf1
    );
  blk00000001_blk0000078d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e2,
      I1 => blk00000001_sig000003c2,
      I2 => blk00000001_sig000003a2,
      I3 => blk00000001_sig00000382,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cf0
    );
  blk00000001_blk0000078c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e3,
      I1 => blk00000001_sig000003c3,
      I2 => blk00000001_sig000003a3,
      I3 => blk00000001_sig00000383,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cef
    );
  blk00000001_blk0000078b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e4,
      I1 => blk00000001_sig000003c4,
      I2 => blk00000001_sig000003a4,
      I3 => blk00000001_sig00000384,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cee
    );
  blk00000001_blk0000078a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e5,
      I1 => blk00000001_sig000003c5,
      I2 => blk00000001_sig000003a5,
      I3 => blk00000001_sig00000385,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ced
    );
  blk00000001_blk00000789 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e6,
      I1 => blk00000001_sig000003c6,
      I2 => blk00000001_sig000003a6,
      I3 => blk00000001_sig00000386,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000cec
    );
  blk00000001_blk00000788 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e7,
      I1 => blk00000001_sig000003c7,
      I2 => blk00000001_sig000003a7,
      I3 => blk00000001_sig00000387,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ceb
    );
  blk00000001_blk00000787 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cfa,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000347
    );
  blk00000001_blk00000786 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000348
    );
  blk00000001_blk00000785 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000349
    );
  blk00000001_blk00000784 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034a
    );
  blk00000001_blk00000783 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034b
    );
  blk00000001_blk00000782 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034c
    );
  blk00000001_blk00000781 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034d
    );
  blk00000001_blk00000780 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034e
    );
  blk00000001_blk0000077f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000034f
    );
  blk00000001_blk0000077e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000350
    );
  blk00000001_blk0000077d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cf0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000351
    );
  blk00000001_blk0000077c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cef,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000352
    );
  blk00000001_blk0000077b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cee,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000353
    );
  blk00000001_blk0000077a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ced,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000354
    );
  blk00000001_blk00000779 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cec,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000355
    );
  blk00000001_blk00000778 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ceb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000356
    );
  blk00000001_blk00000777 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d8,
      I1 => blk00000001_sig000003b8,
      I2 => blk00000001_sig00000398,
      I3 => blk00000001_sig00000378,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cea
    );
  blk00000001_blk00000776 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d9,
      I1 => blk00000001_sig000003b9,
      I2 => blk00000001_sig00000399,
      I3 => blk00000001_sig00000379,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce9
    );
  blk00000001_blk00000775 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003da,
      I1 => blk00000001_sig000003ba,
      I2 => blk00000001_sig0000039a,
      I3 => blk00000001_sig0000037a,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce8
    );
  blk00000001_blk00000774 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003db,
      I1 => blk00000001_sig000003bb,
      I2 => blk00000001_sig0000039b,
      I3 => blk00000001_sig0000037b,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce7
    );
  blk00000001_blk00000773 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dc,
      I1 => blk00000001_sig000003bc,
      I2 => blk00000001_sig0000039c,
      I3 => blk00000001_sig0000037c,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce6
    );
  blk00000001_blk00000772 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003dd,
      I1 => blk00000001_sig000003bd,
      I2 => blk00000001_sig0000039d,
      I3 => blk00000001_sig0000037d,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce5
    );
  blk00000001_blk00000771 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003de,
      I1 => blk00000001_sig000003be,
      I2 => blk00000001_sig0000039e,
      I3 => blk00000001_sig0000037e,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce4
    );
  blk00000001_blk00000770 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003df,
      I1 => blk00000001_sig000003bf,
      I2 => blk00000001_sig0000039f,
      I3 => blk00000001_sig0000037f,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce3
    );
  blk00000001_blk0000076f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e0,
      I1 => blk00000001_sig000003c0,
      I2 => blk00000001_sig000003a0,
      I3 => blk00000001_sig00000380,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce2
    );
  blk00000001_blk0000076e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e1,
      I1 => blk00000001_sig000003c1,
      I2 => blk00000001_sig000003a1,
      I3 => blk00000001_sig00000381,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce1
    );
  blk00000001_blk0000076d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e2,
      I1 => blk00000001_sig000003c2,
      I2 => blk00000001_sig000003a2,
      I3 => blk00000001_sig00000382,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000ce0
    );
  blk00000001_blk0000076c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e3,
      I1 => blk00000001_sig000003c3,
      I2 => blk00000001_sig000003a3,
      I3 => blk00000001_sig00000383,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cdf
    );
  blk00000001_blk0000076b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e4,
      I1 => blk00000001_sig000003c4,
      I2 => blk00000001_sig000003a4,
      I3 => blk00000001_sig00000384,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cde
    );
  blk00000001_blk0000076a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e5,
      I1 => blk00000001_sig000003c5,
      I2 => blk00000001_sig000003a5,
      I3 => blk00000001_sig00000385,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cdd
    );
  blk00000001_blk00000769 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e6,
      I1 => blk00000001_sig000003c6,
      I2 => blk00000001_sig000003a6,
      I3 => blk00000001_sig00000386,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cdc
    );
  blk00000001_blk00000768 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003e7,
      I1 => blk00000001_sig000003c7,
      I2 => blk00000001_sig000003a7,
      I3 => blk00000001_sig00000387,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000cdb
    );
  blk00000001_blk00000767 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cea,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000357
    );
  blk00000001_blk00000766 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000358
    );
  blk00000001_blk00000765 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000359
    );
  blk00000001_blk00000764 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035a
    );
  blk00000001_blk00000763 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035b
    );
  blk00000001_blk00000762 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035c
    );
  blk00000001_blk00000761 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035d
    );
  blk00000001_blk00000760 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035e
    );
  blk00000001_blk0000075f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000035f
    );
  blk00000001_blk0000075e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000360
    );
  blk00000001_blk0000075d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ce0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000361
    );
  blk00000001_blk0000075c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cdf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000362
    );
  blk00000001_blk0000075b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cde,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000363
    );
  blk00000001_blk0000075a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cdd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000364
    );
  blk00000001_blk00000759 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cdc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000365
    );
  blk00000001_blk00000758 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cdb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000366
    );
  blk00000001_blk00000757 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cd1,
      Q => blk00000001_sig00000cd9
    );
  blk00000001_blk00000756 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ccd,
      Q => blk00000001_sig00000cda
    );
  blk00000001_blk00000755 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ccf,
      Q => blk00000001_sig00000cd7
    );
  blk00000001_blk00000754 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ccb,
      Q => blk00000001_sig00000cd8
    );
  blk00000001_blk00000753 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cd0,
      Q => blk00000001_sig00000cd5
    );
  blk00000001_blk00000752 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ccc,
      Q => blk00000001_sig00000cd6
    );
  blk00000001_blk00000751 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cce,
      Q => blk00000001_sig00000cd3
    );
  blk00000001_blk00000750 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cd2,
      Q => blk00000001_sig00000cd4
    );
  blk00000001_blk0000074f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c8,
      I1 => blk00000001_sig000003a8,
      I2 => blk00000001_sig00000388,
      I3 => blk00000001_sig00000368,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cca
    );
  blk00000001_blk0000074e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c9,
      I1 => blk00000001_sig000003a9,
      I2 => blk00000001_sig00000389,
      I3 => blk00000001_sig00000369,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc9
    );
  blk00000001_blk0000074d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ca,
      I1 => blk00000001_sig000003aa,
      I2 => blk00000001_sig0000038a,
      I3 => blk00000001_sig0000036a,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc8
    );
  blk00000001_blk0000074c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cb,
      I1 => blk00000001_sig000003ab,
      I2 => blk00000001_sig0000038b,
      I3 => blk00000001_sig0000036b,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc7
    );
  blk00000001_blk0000074b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cc,
      I1 => blk00000001_sig000003ac,
      I2 => blk00000001_sig0000038c,
      I3 => blk00000001_sig0000036c,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc6
    );
  blk00000001_blk0000074a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cd,
      I1 => blk00000001_sig000003ad,
      I2 => blk00000001_sig0000038d,
      I3 => blk00000001_sig0000036d,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc5
    );
  blk00000001_blk00000749 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ce,
      I1 => blk00000001_sig000003ae,
      I2 => blk00000001_sig0000038e,
      I3 => blk00000001_sig0000036e,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc4
    );
  blk00000001_blk00000748 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cf,
      I1 => blk00000001_sig000003af,
      I2 => blk00000001_sig0000038f,
      I3 => blk00000001_sig0000036f,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc3
    );
  blk00000001_blk00000747 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d0,
      I1 => blk00000001_sig000003b0,
      I2 => blk00000001_sig00000390,
      I3 => blk00000001_sig00000370,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc2
    );
  blk00000001_blk00000746 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d1,
      I1 => blk00000001_sig000003b1,
      I2 => blk00000001_sig00000391,
      I3 => blk00000001_sig00000371,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc1
    );
  blk00000001_blk00000745 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d2,
      I1 => blk00000001_sig000003b2,
      I2 => blk00000001_sig00000392,
      I3 => blk00000001_sig00000372,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cc0
    );
  blk00000001_blk00000744 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d3,
      I1 => blk00000001_sig000003b3,
      I2 => blk00000001_sig00000393,
      I3 => blk00000001_sig00000373,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cbf
    );
  blk00000001_blk00000743 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d4,
      I1 => blk00000001_sig000003b4,
      I2 => blk00000001_sig00000394,
      I3 => blk00000001_sig00000374,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cbe
    );
  blk00000001_blk00000742 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d5,
      I1 => blk00000001_sig000003b5,
      I2 => blk00000001_sig00000395,
      I3 => blk00000001_sig00000375,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cbd
    );
  blk00000001_blk00000741 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d6,
      I1 => blk00000001_sig000003b6,
      I2 => blk00000001_sig00000396,
      I3 => blk00000001_sig00000376,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cbc
    );
  blk00000001_blk00000740 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d7,
      I1 => blk00000001_sig000003b7,
      I2 => blk00000001_sig00000397,
      I3 => blk00000001_sig00000377,
      I4 => blk00000001_sig00000cd5,
      I5 => blk00000001_sig00000cd6,
      O => blk00000001_sig00000cbb
    );
  blk00000001_blk0000073f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cca,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e7
    );
  blk00000001_blk0000073e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e8
    );
  blk00000001_blk0000073d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002e9
    );
  blk00000001_blk0000073c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ea
    );
  blk00000001_blk0000073b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002eb
    );
  blk00000001_blk0000073a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ec
    );
  blk00000001_blk00000739 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ed
    );
  blk00000001_blk00000738 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ee
    );
  blk00000001_blk00000737 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ef
    );
  blk00000001_blk00000736 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f0
    );
  blk00000001_blk00000735 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cc0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f1
    );
  blk00000001_blk00000734 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cbf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f2
    );
  blk00000001_blk00000733 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cbe,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f3
    );
  blk00000001_blk00000732 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cbd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f4
    );
  blk00000001_blk00000731 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cbc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f5
    );
  blk00000001_blk00000730 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cbb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f6
    );
  blk00000001_blk0000072f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c8,
      I1 => blk00000001_sig000003a8,
      I2 => blk00000001_sig00000388,
      I3 => blk00000001_sig00000368,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cba
    );
  blk00000001_blk0000072e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c9,
      I1 => blk00000001_sig000003a9,
      I2 => blk00000001_sig00000389,
      I3 => blk00000001_sig00000369,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb9
    );
  blk00000001_blk0000072d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ca,
      I1 => blk00000001_sig000003aa,
      I2 => blk00000001_sig0000038a,
      I3 => blk00000001_sig0000036a,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb8
    );
  blk00000001_blk0000072c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cb,
      I1 => blk00000001_sig000003ab,
      I2 => blk00000001_sig0000038b,
      I3 => blk00000001_sig0000036b,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb7
    );
  blk00000001_blk0000072b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cc,
      I1 => blk00000001_sig000003ac,
      I2 => blk00000001_sig0000038c,
      I3 => blk00000001_sig0000036c,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb6
    );
  blk00000001_blk0000072a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cd,
      I1 => blk00000001_sig000003ad,
      I2 => blk00000001_sig0000038d,
      I3 => blk00000001_sig0000036d,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb5
    );
  blk00000001_blk00000729 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ce,
      I1 => blk00000001_sig000003ae,
      I2 => blk00000001_sig0000038e,
      I3 => blk00000001_sig0000036e,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb4
    );
  blk00000001_blk00000728 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cf,
      I1 => blk00000001_sig000003af,
      I2 => blk00000001_sig0000038f,
      I3 => blk00000001_sig0000036f,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb3
    );
  blk00000001_blk00000727 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d0,
      I1 => blk00000001_sig000003b0,
      I2 => blk00000001_sig00000390,
      I3 => blk00000001_sig00000370,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb2
    );
  blk00000001_blk00000726 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d1,
      I1 => blk00000001_sig000003b1,
      I2 => blk00000001_sig00000391,
      I3 => blk00000001_sig00000371,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb1
    );
  blk00000001_blk00000725 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d2,
      I1 => blk00000001_sig000003b2,
      I2 => blk00000001_sig00000392,
      I3 => blk00000001_sig00000372,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cb0
    );
  blk00000001_blk00000724 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d3,
      I1 => blk00000001_sig000003b3,
      I2 => blk00000001_sig00000393,
      I3 => blk00000001_sig00000373,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000caf
    );
  blk00000001_blk00000723 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d4,
      I1 => blk00000001_sig000003b4,
      I2 => blk00000001_sig00000394,
      I3 => blk00000001_sig00000374,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cae
    );
  blk00000001_blk00000722 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d5,
      I1 => blk00000001_sig000003b5,
      I2 => blk00000001_sig00000395,
      I3 => blk00000001_sig00000375,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cad
    );
  blk00000001_blk00000721 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d6,
      I1 => blk00000001_sig000003b6,
      I2 => blk00000001_sig00000396,
      I3 => blk00000001_sig00000376,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cac
    );
  blk00000001_blk00000720 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d7,
      I1 => blk00000001_sig000003b7,
      I2 => blk00000001_sig00000397,
      I3 => blk00000001_sig00000377,
      I4 => blk00000001_sig00000cd7,
      I5 => blk00000001_sig00000cd8,
      O => blk00000001_sig00000cab
    );
  blk00000001_blk0000071f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cba,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f7
    );
  blk00000001_blk0000071e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f8
    );
  blk00000001_blk0000071d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002f9
    );
  blk00000001_blk0000071c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002fa
    );
  blk00000001_blk0000071b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002fb
    );
  blk00000001_blk0000071a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002fc
    );
  blk00000001_blk00000719 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002fd
    );
  blk00000001_blk00000718 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002fe
    );
  blk00000001_blk00000717 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000002ff
    );
  blk00000001_blk00000716 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000300
    );
  blk00000001_blk00000715 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cb0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000301
    );
  blk00000001_blk00000714 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000caf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000302
    );
  blk00000001_blk00000713 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cae,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000303
    );
  blk00000001_blk00000712 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cad,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000304
    );
  blk00000001_blk00000711 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cac,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000305
    );
  blk00000001_blk00000710 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000cab,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000306
    );
  blk00000001_blk0000070f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c8,
      I1 => blk00000001_sig000003a8,
      I2 => blk00000001_sig00000388,
      I3 => blk00000001_sig00000368,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000caa
    );
  blk00000001_blk0000070e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c9,
      I1 => blk00000001_sig000003a9,
      I2 => blk00000001_sig00000389,
      I3 => blk00000001_sig00000369,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca9
    );
  blk00000001_blk0000070d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ca,
      I1 => blk00000001_sig000003aa,
      I2 => blk00000001_sig0000038a,
      I3 => blk00000001_sig0000036a,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca8
    );
  blk00000001_blk0000070c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cb,
      I1 => blk00000001_sig000003ab,
      I2 => blk00000001_sig0000038b,
      I3 => blk00000001_sig0000036b,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca7
    );
  blk00000001_blk0000070b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cc,
      I1 => blk00000001_sig000003ac,
      I2 => blk00000001_sig0000038c,
      I3 => blk00000001_sig0000036c,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca6
    );
  blk00000001_blk0000070a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cd,
      I1 => blk00000001_sig000003ad,
      I2 => blk00000001_sig0000038d,
      I3 => blk00000001_sig0000036d,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca5
    );
  blk00000001_blk00000709 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ce,
      I1 => blk00000001_sig000003ae,
      I2 => blk00000001_sig0000038e,
      I3 => blk00000001_sig0000036e,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca4
    );
  blk00000001_blk00000708 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cf,
      I1 => blk00000001_sig000003af,
      I2 => blk00000001_sig0000038f,
      I3 => blk00000001_sig0000036f,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca3
    );
  blk00000001_blk00000707 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d0,
      I1 => blk00000001_sig000003b0,
      I2 => blk00000001_sig00000390,
      I3 => blk00000001_sig00000370,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca2
    );
  blk00000001_blk00000706 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d1,
      I1 => blk00000001_sig000003b1,
      I2 => blk00000001_sig00000391,
      I3 => blk00000001_sig00000371,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca1
    );
  blk00000001_blk00000705 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d2,
      I1 => blk00000001_sig000003b2,
      I2 => blk00000001_sig00000392,
      I3 => blk00000001_sig00000372,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000ca0
    );
  blk00000001_blk00000704 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d3,
      I1 => blk00000001_sig000003b3,
      I2 => blk00000001_sig00000393,
      I3 => blk00000001_sig00000373,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000c9f
    );
  blk00000001_blk00000703 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d4,
      I1 => blk00000001_sig000003b4,
      I2 => blk00000001_sig00000394,
      I3 => blk00000001_sig00000374,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000c9e
    );
  blk00000001_blk00000702 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d5,
      I1 => blk00000001_sig000003b5,
      I2 => blk00000001_sig00000395,
      I3 => blk00000001_sig00000375,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000c9d
    );
  blk00000001_blk00000701 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d6,
      I1 => blk00000001_sig000003b6,
      I2 => blk00000001_sig00000396,
      I3 => blk00000001_sig00000376,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000c9c
    );
  blk00000001_blk00000700 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d7,
      I1 => blk00000001_sig000003b7,
      I2 => blk00000001_sig00000397,
      I3 => blk00000001_sig00000377,
      I4 => blk00000001_sig00000cd9,
      I5 => blk00000001_sig00000cda,
      O => blk00000001_sig00000c9b
    );
  blk00000001_blk000006ff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000caa,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000307
    );
  blk00000001_blk000006fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000308
    );
  blk00000001_blk000006fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000309
    );
  blk00000001_blk000006fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030a
    );
  blk00000001_blk000006fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030b
    );
  blk00000001_blk000006fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030c
    );
  blk00000001_blk000006f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030d
    );
  blk00000001_blk000006f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030e
    );
  blk00000001_blk000006f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000030f
    );
  blk00000001_blk000006f6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000310
    );
  blk00000001_blk000006f5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000ca0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000311
    );
  blk00000001_blk000006f4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000312
    );
  blk00000001_blk000006f3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000313
    );
  blk00000001_blk000006f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000314
    );
  blk00000001_blk000006f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000315
    );
  blk00000001_blk000006f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000316
    );
  blk00000001_blk000006ef : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c8,
      I1 => blk00000001_sig000003a8,
      I2 => blk00000001_sig00000388,
      I3 => blk00000001_sig00000368,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c9a
    );
  blk00000001_blk000006ee : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003c9,
      I1 => blk00000001_sig000003a9,
      I2 => blk00000001_sig00000389,
      I3 => blk00000001_sig00000369,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c99
    );
  blk00000001_blk000006ed : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ca,
      I1 => blk00000001_sig000003aa,
      I2 => blk00000001_sig0000038a,
      I3 => blk00000001_sig0000036a,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c98
    );
  blk00000001_blk000006ec : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cb,
      I1 => blk00000001_sig000003ab,
      I2 => blk00000001_sig0000038b,
      I3 => blk00000001_sig0000036b,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c97
    );
  blk00000001_blk000006eb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cc,
      I1 => blk00000001_sig000003ac,
      I2 => blk00000001_sig0000038c,
      I3 => blk00000001_sig0000036c,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c96
    );
  blk00000001_blk000006ea : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cd,
      I1 => blk00000001_sig000003ad,
      I2 => blk00000001_sig0000038d,
      I3 => blk00000001_sig0000036d,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c95
    );
  blk00000001_blk000006e9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003ce,
      I1 => blk00000001_sig000003ae,
      I2 => blk00000001_sig0000038e,
      I3 => blk00000001_sig0000036e,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c94
    );
  blk00000001_blk000006e8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003cf,
      I1 => blk00000001_sig000003af,
      I2 => blk00000001_sig0000038f,
      I3 => blk00000001_sig0000036f,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c93
    );
  blk00000001_blk000006e7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d0,
      I1 => blk00000001_sig000003b0,
      I2 => blk00000001_sig00000390,
      I3 => blk00000001_sig00000370,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c92
    );
  blk00000001_blk000006e6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d1,
      I1 => blk00000001_sig000003b1,
      I2 => blk00000001_sig00000391,
      I3 => blk00000001_sig00000371,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c91
    );
  blk00000001_blk000006e5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d2,
      I1 => blk00000001_sig000003b2,
      I2 => blk00000001_sig00000392,
      I3 => blk00000001_sig00000372,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c90
    );
  blk00000001_blk000006e4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d3,
      I1 => blk00000001_sig000003b3,
      I2 => blk00000001_sig00000393,
      I3 => blk00000001_sig00000373,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c8f
    );
  blk00000001_blk000006e3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d4,
      I1 => blk00000001_sig000003b4,
      I2 => blk00000001_sig00000394,
      I3 => blk00000001_sig00000374,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c8e
    );
  blk00000001_blk000006e2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d5,
      I1 => blk00000001_sig000003b5,
      I2 => blk00000001_sig00000395,
      I3 => blk00000001_sig00000375,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c8d
    );
  blk00000001_blk000006e1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d6,
      I1 => blk00000001_sig000003b6,
      I2 => blk00000001_sig00000396,
      I3 => blk00000001_sig00000376,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c8c
    );
  blk00000001_blk000006e0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000003d7,
      I1 => blk00000001_sig000003b7,
      I2 => blk00000001_sig00000397,
      I3 => blk00000001_sig00000377,
      I4 => blk00000001_sig00000cd3,
      I5 => blk00000001_sig00000cd4,
      O => blk00000001_sig00000c8b
    );
  blk00000001_blk000006df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c9a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000317
    );
  blk00000001_blk000006de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c99,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000318
    );
  blk00000001_blk000006dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c98,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000319
    );
  blk00000001_blk000006dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c97,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031a
    );
  blk00000001_blk000006db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c96,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031b
    );
  blk00000001_blk000006da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c95,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031c
    );
  blk00000001_blk000006d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c94,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031d
    );
  blk00000001_blk000006d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c93,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031e
    );
  blk00000001_blk000006d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c92,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000031f
    );
  blk00000001_blk000006d6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c91,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000320
    );
  blk00000001_blk000006d5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c90,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000321
    );
  blk00000001_blk000006d4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000322
    );
  blk00000001_blk000006d3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000323
    );
  blk00000001_blk000006d2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000324
    );
  blk00000001_blk000006d1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000325
    );
  blk00000001_blk000006d0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000326
    );
  blk00000001_blk000006cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000c8a,
      Q => blk00000001_sig00000367
    );
  blk00000001_blk000006ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001ad,
      Q => blk00000001_sig00000ba0
    );
  blk00000001_blk000006cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001ad,
      Q => blk00000001_sig00000b9e
    );
  blk00000001_blk000006cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5f,
      Q => blk00000001_sig00000acc
    );
  blk00000001_blk000006cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b60,
      Q => blk00000001_sig00000acd
    );
  blk00000001_blk000006ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b61,
      Q => blk00000001_sig00000ace
    );
  blk00000001_blk000006c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b62,
      Q => blk00000001_sig00000acf
    );
  blk00000001_blk000006c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b63,
      Q => blk00000001_sig00000ad0
    );
  blk00000001_blk000006c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b64,
      Q => blk00000001_sig00000ad1
    );
  blk00000001_blk000006c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b65,
      Q => blk00000001_sig00000ad2
    );
  blk00000001_blk000006c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b66,
      Q => blk00000001_sig00000ad3
    );
  blk00000001_blk000006c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b67,
      Q => blk00000001_sig00000ad4
    );
  blk00000001_blk000006c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b68,
      Q => blk00000001_sig00000ad5
    );
  blk00000001_blk000006c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b69,
      Q => blk00000001_sig00000ad6
    );
  blk00000001_blk000006c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6a,
      Q => blk00000001_sig00000ad7
    );
  blk00000001_blk000006c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6b,
      Q => blk00000001_sig00000ad8
    );
  blk00000001_blk000006bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6c,
      Q => blk00000001_sig00000ad9
    );
  blk00000001_blk000006be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6d,
      Q => blk00000001_sig00000ada
    );
  blk00000001_blk000006bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6e,
      Q => blk00000001_sig00000adb
    );
  blk00000001_blk000006bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b6f,
      Q => blk00000001_sig00000adc
    );
  blk00000001_blk000006bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b70,
      Q => blk00000001_sig00000add
    );
  blk00000001_blk000006ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b71,
      Q => blk00000001_sig00000ade
    );
  blk00000001_blk000006b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b72,
      Q => blk00000001_sig00000adf
    );
  blk00000001_blk000006b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b73,
      Q => blk00000001_sig00000ae0
    );
  blk00000001_blk000006b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b74,
      Q => blk00000001_sig00000ae1
    );
  blk00000001_blk000006b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b75,
      Q => blk00000001_sig00000ae2
    );
  blk00000001_blk000006b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b76,
      Q => blk00000001_sig00000ae3
    );
  blk00000001_blk000006b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b77,
      Q => blk00000001_sig00000ae4
    );
  blk00000001_blk000006b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b78,
      Q => blk00000001_sig00000ae5
    );
  blk00000001_blk000006b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b79,
      Q => blk00000001_sig00000ae6
    );
  blk00000001_blk000006b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7a,
      Q => blk00000001_sig00000ae7
    );
  blk00000001_blk000006b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7b,
      Q => blk00000001_sig00000ae8
    );
  blk00000001_blk000006af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7c,
      Q => blk00000001_sig00000ae9
    );
  blk00000001_blk000006ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7d,
      Q => blk00000001_sig00000aea
    );
  blk00000001_blk000006ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7e,
      Q => blk00000001_sig00000aeb
    );
  blk00000001_blk000006ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b7f,
      Q => blk00000001_sig00000aec
    );
  blk00000001_blk000006ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b80,
      Q => blk00000001_sig00000aed
    );
  blk00000001_blk000006aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b81,
      Q => blk00000001_sig00000aee
    );
  blk00000001_blk000006a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b82,
      Q => blk00000001_sig00000aef
    );
  blk00000001_blk000006a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b83,
      Q => blk00000001_sig00000af0
    );
  blk00000001_blk000006a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b84,
      Q => blk00000001_sig00000af1
    );
  blk00000001_blk000006a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b85,
      Q => blk00000001_sig00000af2
    );
  blk00000001_blk000006a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b86,
      Q => blk00000001_sig00000af3
    );
  blk00000001_blk000006a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b87,
      Q => blk00000001_sig00000af4
    );
  blk00000001_blk000006a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b88,
      Q => blk00000001_sig00000af5
    );
  blk00000001_blk000006a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4a,
      Q => blk00000001_sig00000ab7
    );
  blk00000001_blk000006a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4b,
      Q => blk00000001_sig00000ab8
    );
  blk00000001_blk000006a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4c,
      Q => blk00000001_sig00000ab9
    );
  blk00000001_blk0000069f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4d,
      Q => blk00000001_sig00000aba
    );
  blk00000001_blk0000069e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4e,
      Q => blk00000001_sig00000abb
    );
  blk00000001_blk0000069d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b4f,
      Q => blk00000001_sig00000abc
    );
  blk00000001_blk0000069c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b50,
      Q => blk00000001_sig00000abd
    );
  blk00000001_blk0000069b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b51,
      Q => blk00000001_sig00000abe
    );
  blk00000001_blk0000069a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b52,
      Q => blk00000001_sig00000abf
    );
  blk00000001_blk00000699 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b53,
      Q => blk00000001_sig00000ac0
    );
  blk00000001_blk00000698 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b54,
      Q => blk00000001_sig00000ac1
    );
  blk00000001_blk00000697 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b55,
      Q => blk00000001_sig00000ac2
    );
  blk00000001_blk00000696 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b56,
      Q => blk00000001_sig00000ac3
    );
  blk00000001_blk00000695 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b57,
      Q => blk00000001_sig00000ac4
    );
  blk00000001_blk00000694 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b58,
      Q => blk00000001_sig00000ac5
    );
  blk00000001_blk00000693 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b59,
      Q => blk00000001_sig00000ac6
    );
  blk00000001_blk00000692 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5a,
      Q => blk00000001_sig00000ac7
    );
  blk00000001_blk00000691 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5b,
      Q => blk00000001_sig00000ac8
    );
  blk00000001_blk00000690 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5c,
      Q => blk00000001_sig00000ac9
    );
  blk00000001_blk0000068f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5d,
      Q => blk00000001_sig00000aca
    );
  blk00000001_blk0000068e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b5e,
      Q => blk00000001_sig00000acb
    );
  blk00000001_blk0000068d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b89,
      Q => blk00000001_sig00000a4e
    );
  blk00000001_blk0000068c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8a,
      Q => blk00000001_sig00000a4f
    );
  blk00000001_blk0000068b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8b,
      Q => blk00000001_sig00000a50
    );
  blk00000001_blk0000068a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8c,
      Q => blk00000001_sig00000a51
    );
  blk00000001_blk00000689 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8d,
      Q => blk00000001_sig00000a52
    );
  blk00000001_blk00000688 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8e,
      Q => blk00000001_sig00000a53
    );
  blk00000001_blk00000687 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b8f,
      Q => blk00000001_sig00000a54
    );
  blk00000001_blk00000686 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b90,
      Q => blk00000001_sig00000a55
    );
  blk00000001_blk00000685 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b91,
      Q => blk00000001_sig00000a56
    );
  blk00000001_blk00000684 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b92,
      Q => blk00000001_sig00000a57
    );
  blk00000001_blk00000683 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b93,
      Q => blk00000001_sig00000a58
    );
  blk00000001_blk00000682 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b94,
      Q => blk00000001_sig00000a59
    );
  blk00000001_blk00000681 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b95,
      Q => blk00000001_sig00000a5a
    );
  blk00000001_blk00000680 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b96,
      Q => blk00000001_sig00000a5b
    );
  blk00000001_blk0000067f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b97,
      Q => blk00000001_sig00000a5c
    );
  blk00000001_blk0000067e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b98,
      Q => blk00000001_sig00000a5d
    );
  blk00000001_blk0000067d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b99,
      Q => blk00000001_sig00000a5e
    );
  blk00000001_blk0000067c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b9a,
      Q => blk00000001_sig00000a5f
    );
  blk00000001_blk0000067b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b9b,
      Q => blk00000001_sig00000a60
    );
  blk00000001_blk0000067a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b9c,
      Q => blk00000001_sig00000a61
    );
  blk00000001_blk00000679 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b9d,
      Q => blk00000001_sig00000a62
    );
  blk00000001_blk00000678 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b20,
      Q => blk00000001_sig00000a8d
    );
  blk00000001_blk00000677 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b21,
      Q => blk00000001_sig00000a8e
    );
  blk00000001_blk00000676 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b22,
      Q => blk00000001_sig00000a8f
    );
  blk00000001_blk00000675 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b23,
      Q => blk00000001_sig00000a90
    );
  blk00000001_blk00000674 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b24,
      Q => blk00000001_sig00000a91
    );
  blk00000001_blk00000673 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b25,
      Q => blk00000001_sig00000a92
    );
  blk00000001_blk00000672 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b26,
      Q => blk00000001_sig00000a93
    );
  blk00000001_blk00000671 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b27,
      Q => blk00000001_sig00000a94
    );
  blk00000001_blk00000670 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b28,
      Q => blk00000001_sig00000a95
    );
  blk00000001_blk0000066f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b29,
      Q => blk00000001_sig00000a96
    );
  blk00000001_blk0000066e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2a,
      Q => blk00000001_sig00000a97
    );
  blk00000001_blk0000066d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2b,
      Q => blk00000001_sig00000a98
    );
  blk00000001_blk0000066c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2c,
      Q => blk00000001_sig00000a99
    );
  blk00000001_blk0000066b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2d,
      Q => blk00000001_sig00000a9a
    );
  blk00000001_blk0000066a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2e,
      Q => blk00000001_sig00000a9b
    );
  blk00000001_blk00000669 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b2f,
      Q => blk00000001_sig00000a9c
    );
  blk00000001_blk00000668 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b30,
      Q => blk00000001_sig00000a9d
    );
  blk00000001_blk00000667 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b31,
      Q => blk00000001_sig00000a9e
    );
  blk00000001_blk00000666 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b32,
      Q => blk00000001_sig00000a9f
    );
  blk00000001_blk00000665 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b33,
      Q => blk00000001_sig00000aa0
    );
  blk00000001_blk00000664 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b34,
      Q => blk00000001_sig00000aa1
    );
  blk00000001_blk00000663 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b35,
      Q => blk00000001_sig00000aa2
    );
  blk00000001_blk00000662 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b36,
      Q => blk00000001_sig00000aa3
    );
  blk00000001_blk00000661 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b37,
      Q => blk00000001_sig00000aa4
    );
  blk00000001_blk00000660 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b38,
      Q => blk00000001_sig00000aa5
    );
  blk00000001_blk0000065f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b39,
      Q => blk00000001_sig00000aa6
    );
  blk00000001_blk0000065e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3a,
      Q => blk00000001_sig00000aa7
    );
  blk00000001_blk0000065d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3b,
      Q => blk00000001_sig00000aa8
    );
  blk00000001_blk0000065c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3c,
      Q => blk00000001_sig00000aa9
    );
  blk00000001_blk0000065b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3d,
      Q => blk00000001_sig00000aaa
    );
  blk00000001_blk0000065a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3e,
      Q => blk00000001_sig00000aab
    );
  blk00000001_blk00000659 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b3f,
      Q => blk00000001_sig00000aac
    );
  blk00000001_blk00000658 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b40,
      Q => blk00000001_sig00000aad
    );
  blk00000001_blk00000657 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b41,
      Q => blk00000001_sig00000aae
    );
  blk00000001_blk00000656 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b42,
      Q => blk00000001_sig00000aaf
    );
  blk00000001_blk00000655 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b43,
      Q => blk00000001_sig00000ab0
    );
  blk00000001_blk00000654 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b44,
      Q => blk00000001_sig00000ab1
    );
  blk00000001_blk00000653 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b45,
      Q => blk00000001_sig00000ab2
    );
  blk00000001_blk00000652 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b46,
      Q => blk00000001_sig00000ab3
    );
  blk00000001_blk00000651 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b47,
      Q => blk00000001_sig00000ab4
    );
  blk00000001_blk00000650 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b48,
      Q => blk00000001_sig00000ab5
    );
  blk00000001_blk0000064f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b49,
      Q => blk00000001_sig00000ab6
    );
  blk00000001_blk0000064e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0b,
      Q => blk00000001_sig00000a78
    );
  blk00000001_blk0000064d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0c,
      Q => blk00000001_sig00000a79
    );
  blk00000001_blk0000064c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0d,
      Q => blk00000001_sig00000a7a
    );
  blk00000001_blk0000064b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0e,
      Q => blk00000001_sig00000a7b
    );
  blk00000001_blk0000064a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0f,
      Q => blk00000001_sig00000a7c
    );
  blk00000001_blk00000649 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b10,
      Q => blk00000001_sig00000a7d
    );
  blk00000001_blk00000648 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b11,
      Q => blk00000001_sig00000a7e
    );
  blk00000001_blk00000647 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b12,
      Q => blk00000001_sig00000a7f
    );
  blk00000001_blk00000646 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b13,
      Q => blk00000001_sig00000a80
    );
  blk00000001_blk00000645 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b14,
      Q => blk00000001_sig00000a81
    );
  blk00000001_blk00000644 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b15,
      Q => blk00000001_sig00000a82
    );
  blk00000001_blk00000643 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b16,
      Q => blk00000001_sig00000a83
    );
  blk00000001_blk00000642 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b17,
      Q => blk00000001_sig00000a84
    );
  blk00000001_blk00000641 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b18,
      Q => blk00000001_sig00000a85
    );
  blk00000001_blk00000640 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b19,
      Q => blk00000001_sig00000a86
    );
  blk00000001_blk0000063f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1a,
      Q => blk00000001_sig00000a87
    );
  blk00000001_blk0000063e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1b,
      Q => blk00000001_sig00000a88
    );
  blk00000001_blk0000063d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1c,
      Q => blk00000001_sig00000a89
    );
  blk00000001_blk0000063c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1d,
      Q => blk00000001_sig00000a8a
    );
  blk00000001_blk0000063b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1e,
      Q => blk00000001_sig00000a8b
    );
  blk00000001_blk0000063a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b1f,
      Q => blk00000001_sig00000a8c
    );
  blk00000001_blk00000639 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000af6,
      Q => blk00000001_sig00000a63
    );
  blk00000001_blk00000638 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000af7,
      Q => blk00000001_sig00000a64
    );
  blk00000001_blk00000637 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000af8,
      Q => blk00000001_sig00000a65
    );
  blk00000001_blk00000636 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000af9,
      Q => blk00000001_sig00000a66
    );
  blk00000001_blk00000635 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000afa,
      Q => blk00000001_sig00000a67
    );
  blk00000001_blk00000634 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000afb,
      Q => blk00000001_sig00000a68
    );
  blk00000001_blk00000633 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000afc,
      Q => blk00000001_sig00000a69
    );
  blk00000001_blk00000632 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000afd,
      Q => blk00000001_sig00000a6a
    );
  blk00000001_blk00000631 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000afe,
      Q => blk00000001_sig00000a6b
    );
  blk00000001_blk00000630 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000aff,
      Q => blk00000001_sig00000a6c
    );
  blk00000001_blk0000062f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b00,
      Q => blk00000001_sig00000a6d
    );
  blk00000001_blk0000062e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b01,
      Q => blk00000001_sig00000a6e
    );
  blk00000001_blk0000062d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b02,
      Q => blk00000001_sig00000a6f
    );
  blk00000001_blk0000062c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b03,
      Q => blk00000001_sig00000a70
    );
  blk00000001_blk0000062b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b04,
      Q => blk00000001_sig00000a71
    );
  blk00000001_blk0000062a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b05,
      Q => blk00000001_sig00000a72
    );
  blk00000001_blk00000629 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b06,
      Q => blk00000001_sig00000a73
    );
  blk00000001_blk00000628 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b07,
      Q => blk00000001_sig00000a74
    );
  blk00000001_blk00000627 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b08,
      Q => blk00000001_sig00000a75
    );
  blk00000001_blk00000626 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b09,
      Q => blk00000001_sig00000a76
    );
  blk00000001_blk00000625 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000b0a,
      Q => blk00000001_sig00000a77
    );
  blk00000001_blk00000624 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a4d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006c8
    );
  blk00000001_blk00000623 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a4c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006c7
    );
  blk00000001_blk00000622 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a4b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006c6
    );
  blk00000001_blk00000621 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a4a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000377
    );
  blk00000001_blk00000620 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a49,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000376
    );
  blk00000001_blk0000061f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a48,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000375
    );
  blk00000001_blk0000061e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a47,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000374
    );
  blk00000001_blk0000061d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a46,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000373
    );
  blk00000001_blk0000061c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a45,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000372
    );
  blk00000001_blk0000061b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a44,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000371
    );
  blk00000001_blk0000061a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a43,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000370
    );
  blk00000001_blk00000619 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a42,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036f
    );
  blk00000001_blk00000618 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a41,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036e
    );
  blk00000001_blk00000617 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a40,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036d
    );
  blk00000001_blk00000616 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036c
    );
  blk00000001_blk00000615 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036b
    );
  blk00000001_blk00000614 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000036a
    );
  blk00000001_blk00000613 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000369
    );
  blk00000001_blk00000612 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000368
    );
  blk00000001_blk00000611 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a3a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000611_Q_UNCONNECTED
    );
  blk00000001_blk00000610 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a39,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000610_Q_UNCONNECTED
    );
  blk00000001_blk0000060f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a38,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000060f_Q_UNCONNECTED
    );
  blk00000001_blk0000060e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a37,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000060e_Q_UNCONNECTED
    );
  blk00000001_blk0000060d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a36,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000060d_Q_UNCONNECTED
    );
  blk00000001_blk0000060c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a35,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000060c_Q_UNCONNECTED
    );
  blk00000001_blk0000060b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000517,
      I1 => blk00000001_sig00000517,
      I2 => blk00000001_sig00000517,
      I3 => blk00000001_sig00000517,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a4d
    );
  blk00000001_blk0000060a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000516,
      I1 => blk00000001_sig00000517,
      I2 => blk00000001_sig00000517,
      I3 => blk00000001_sig00000517,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a4c
    );
  blk00000001_blk00000609 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000515,
      I1 => blk00000001_sig00000516,
      I2 => blk00000001_sig00000517,
      I3 => blk00000001_sig00000517,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a4b
    );
  blk00000001_blk00000608 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000514,
      I1 => blk00000001_sig00000515,
      I2 => blk00000001_sig00000516,
      I3 => blk00000001_sig00000517,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a4a
    );
  blk00000001_blk00000607 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000513,
      I1 => blk00000001_sig00000514,
      I2 => blk00000001_sig00000515,
      I3 => blk00000001_sig00000516,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a49
    );
  blk00000001_blk00000606 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000512,
      I1 => blk00000001_sig00000513,
      I2 => blk00000001_sig00000514,
      I3 => blk00000001_sig00000515,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a48
    );
  blk00000001_blk00000605 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000511,
      I1 => blk00000001_sig00000512,
      I2 => blk00000001_sig00000513,
      I3 => blk00000001_sig00000514,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a47
    );
  blk00000001_blk00000604 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000510,
      I1 => blk00000001_sig00000511,
      I2 => blk00000001_sig00000512,
      I3 => blk00000001_sig00000513,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a46
    );
  blk00000001_blk00000603 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050f,
      I1 => blk00000001_sig00000510,
      I2 => blk00000001_sig00000511,
      I3 => blk00000001_sig00000512,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a45
    );
  blk00000001_blk00000602 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050e,
      I1 => blk00000001_sig0000050f,
      I2 => blk00000001_sig00000510,
      I3 => blk00000001_sig00000511,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a44
    );
  blk00000001_blk00000601 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050d,
      I1 => blk00000001_sig0000050e,
      I2 => blk00000001_sig0000050f,
      I3 => blk00000001_sig00000510,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a43
    );
  blk00000001_blk00000600 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050c,
      I1 => blk00000001_sig0000050d,
      I2 => blk00000001_sig0000050e,
      I3 => blk00000001_sig0000050f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a42
    );
  blk00000001_blk000005ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050b,
      I1 => blk00000001_sig0000050c,
      I2 => blk00000001_sig0000050d,
      I3 => blk00000001_sig0000050e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a41
    );
  blk00000001_blk000005fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000050a,
      I1 => blk00000001_sig0000050b,
      I2 => blk00000001_sig0000050c,
      I3 => blk00000001_sig0000050d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a40
    );
  blk00000001_blk000005fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000509,
      I1 => blk00000001_sig0000050a,
      I2 => blk00000001_sig0000050b,
      I3 => blk00000001_sig0000050c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3f
    );
  blk00000001_blk000005fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000508,
      I1 => blk00000001_sig00000509,
      I2 => blk00000001_sig0000050a,
      I3 => blk00000001_sig0000050b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3e
    );
  blk00000001_blk000005fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000507,
      I1 => blk00000001_sig00000508,
      I2 => blk00000001_sig00000509,
      I3 => blk00000001_sig0000050a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3d
    );
  blk00000001_blk000005fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000506,
      I1 => blk00000001_sig00000507,
      I2 => blk00000001_sig00000508,
      I3 => blk00000001_sig00000509,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3c
    );
  blk00000001_blk000005f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000505,
      I1 => blk00000001_sig00000506,
      I2 => blk00000001_sig00000507,
      I3 => blk00000001_sig00000508,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3b
    );
  blk00000001_blk000005f8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000504,
      I1 => blk00000001_sig00000505,
      I2 => blk00000001_sig00000506,
      I3 => blk00000001_sig00000507,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a3a
    );
  blk00000001_blk000005f7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000503,
      I1 => blk00000001_sig00000504,
      I2 => blk00000001_sig00000505,
      I3 => blk00000001_sig00000506,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a39
    );
  blk00000001_blk000005f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000502,
      I1 => blk00000001_sig00000503,
      I2 => blk00000001_sig00000504,
      I3 => blk00000001_sig00000505,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a38
    );
  blk00000001_blk000005f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000502,
      I2 => blk00000001_sig00000503,
      I3 => blk00000001_sig00000504,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a37
    );
  blk00000001_blk000005f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000502,
      I3 => blk00000001_sig00000503,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a36
    );
  blk00000001_blk000005f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig00000502,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a35
    );
  blk00000001_blk000005f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a34,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006cb
    );
  blk00000001_blk000005f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a33,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006ca
    );
  blk00000001_blk000005f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a32,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006c9
    );
  blk00000001_blk000005ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a31,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000387
    );
  blk00000001_blk000005ee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a30,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000386
    );
  blk00000001_blk000005ed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000385
    );
  blk00000001_blk000005ec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000384
    );
  blk00000001_blk000005eb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000383
    );
  blk00000001_blk000005ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000382
    );
  blk00000001_blk000005e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000381
    );
  blk00000001_blk000005e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a2a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000380
    );
  blk00000001_blk000005e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a29,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037f
    );
  blk00000001_blk000005e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a28,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037e
    );
  blk00000001_blk000005e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a27,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037d
    );
  blk00000001_blk000005e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a26,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037c
    );
  blk00000001_blk000005e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a25,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037b
    );
  blk00000001_blk000005e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a24,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000037a
    );
  blk00000001_blk000005e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a23,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000379
    );
  blk00000001_blk000005e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a22,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000378
    );
  blk00000001_blk000005df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a21,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005df_Q_UNCONNECTED
    );
  blk00000001_blk000005de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a20,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005de_Q_UNCONNECTED
    );
  blk00000001_blk000005dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005dd_Q_UNCONNECTED
    );
  blk00000001_blk000005dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005dc_Q_UNCONNECTED
    );
  blk00000001_blk000005db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005db_Q_UNCONNECTED
    );
  blk00000001_blk000005da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005da_Q_UNCONNECTED
    );
  blk00000001_blk000005d9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052d,
      I1 => blk00000001_sig0000052d,
      I2 => blk00000001_sig0000052d,
      I3 => blk00000001_sig0000052d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a34
    );
  blk00000001_blk000005d8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052c,
      I1 => blk00000001_sig0000052d,
      I2 => blk00000001_sig0000052d,
      I3 => blk00000001_sig0000052d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a33
    );
  blk00000001_blk000005d7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052b,
      I1 => blk00000001_sig0000052c,
      I2 => blk00000001_sig0000052d,
      I3 => blk00000001_sig0000052d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a32
    );
  blk00000001_blk000005d6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052a,
      I1 => blk00000001_sig0000052b,
      I2 => blk00000001_sig0000052c,
      I3 => blk00000001_sig0000052d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a31
    );
  blk00000001_blk000005d5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000529,
      I1 => blk00000001_sig0000052a,
      I2 => blk00000001_sig0000052b,
      I3 => blk00000001_sig0000052c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a30
    );
  blk00000001_blk000005d4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000528,
      I1 => blk00000001_sig00000529,
      I2 => blk00000001_sig0000052a,
      I3 => blk00000001_sig0000052b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2f
    );
  blk00000001_blk000005d3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000527,
      I1 => blk00000001_sig00000528,
      I2 => blk00000001_sig00000529,
      I3 => blk00000001_sig0000052a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2e
    );
  blk00000001_blk000005d2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000526,
      I1 => blk00000001_sig00000527,
      I2 => blk00000001_sig00000528,
      I3 => blk00000001_sig00000529,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2d
    );
  blk00000001_blk000005d1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000525,
      I1 => blk00000001_sig00000526,
      I2 => blk00000001_sig00000527,
      I3 => blk00000001_sig00000528,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2c
    );
  blk00000001_blk000005d0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000524,
      I1 => blk00000001_sig00000525,
      I2 => blk00000001_sig00000526,
      I3 => blk00000001_sig00000527,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2b
    );
  blk00000001_blk000005cf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000523,
      I1 => blk00000001_sig00000524,
      I2 => blk00000001_sig00000525,
      I3 => blk00000001_sig00000526,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a2a
    );
  blk00000001_blk000005ce : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000522,
      I1 => blk00000001_sig00000523,
      I2 => blk00000001_sig00000524,
      I3 => blk00000001_sig00000525,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a29
    );
  blk00000001_blk000005cd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000521,
      I1 => blk00000001_sig00000522,
      I2 => blk00000001_sig00000523,
      I3 => blk00000001_sig00000524,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a28
    );
  blk00000001_blk000005cc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000520,
      I1 => blk00000001_sig00000521,
      I2 => blk00000001_sig00000522,
      I3 => blk00000001_sig00000523,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a27
    );
  blk00000001_blk000005cb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051f,
      I1 => blk00000001_sig00000520,
      I2 => blk00000001_sig00000521,
      I3 => blk00000001_sig00000522,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a26
    );
  blk00000001_blk000005ca : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051e,
      I1 => blk00000001_sig0000051f,
      I2 => blk00000001_sig00000520,
      I3 => blk00000001_sig00000521,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a25
    );
  blk00000001_blk000005c9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051d,
      I1 => blk00000001_sig0000051e,
      I2 => blk00000001_sig0000051f,
      I3 => blk00000001_sig00000520,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a24
    );
  blk00000001_blk000005c8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051c,
      I1 => blk00000001_sig0000051d,
      I2 => blk00000001_sig0000051e,
      I3 => blk00000001_sig0000051f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a23
    );
  blk00000001_blk000005c7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051b,
      I1 => blk00000001_sig0000051c,
      I2 => blk00000001_sig0000051d,
      I3 => blk00000001_sig0000051e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a22
    );
  blk00000001_blk000005c6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000051a,
      I1 => blk00000001_sig0000051b,
      I2 => blk00000001_sig0000051c,
      I3 => blk00000001_sig0000051d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a21
    );
  blk00000001_blk000005c5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000519,
      I1 => blk00000001_sig0000051a,
      I2 => blk00000001_sig0000051b,
      I3 => blk00000001_sig0000051c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a20
    );
  blk00000001_blk000005c4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000518,
      I1 => blk00000001_sig00000519,
      I2 => blk00000001_sig0000051a,
      I3 => blk00000001_sig0000051b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1f
    );
  blk00000001_blk000005c3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000518,
      I2 => blk00000001_sig00000519,
      I3 => blk00000001_sig0000051a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1e
    );
  blk00000001_blk000005c2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000518,
      I3 => blk00000001_sig00000519,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1d
    );
  blk00000001_blk000005c1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig00000518,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1c
    );
  blk00000001_blk000005c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006ce
    );
  blk00000001_blk000005bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a1a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006cd
    );
  blk00000001_blk000005be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a19,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006cc
    );
  blk00000001_blk000005bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a18,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000397
    );
  blk00000001_blk000005bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a17,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000396
    );
  blk00000001_blk000005bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a16,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000395
    );
  blk00000001_blk000005ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a15,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000394
    );
  blk00000001_blk000005b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a14,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000393
    );
  blk00000001_blk000005b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a13,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000392
    );
  blk00000001_blk000005b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a12,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000391
    );
  blk00000001_blk000005b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a11,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000390
    );
  blk00000001_blk000005b5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a10,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038f
    );
  blk00000001_blk000005b4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038e
    );
  blk00000001_blk000005b3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038d
    );
  blk00000001_blk000005b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038c
    );
  blk00000001_blk000005b1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038b
    );
  blk00000001_blk000005b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000038a
    );
  blk00000001_blk000005af : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a0a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000389
    );
  blk00000001_blk000005ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a09,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000388
    );
  blk00000001_blk000005ad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a08,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005ad_Q_UNCONNECTED
    );
  blk00000001_blk000005ac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a07,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005ac_Q_UNCONNECTED
    );
  blk00000001_blk000005ab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a06,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005ab_Q_UNCONNECTED
    );
  blk00000001_blk000005aa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a05,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005aa_Q_UNCONNECTED
    );
  blk00000001_blk000005a9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a04,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005a9_Q_UNCONNECTED
    );
  blk00000001_blk000005a8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a03,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000005a8_Q_UNCONNECTED
    );
  blk00000001_blk000005a7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000543,
      I1 => blk00000001_sig00000543,
      I2 => blk00000001_sig00000543,
      I3 => blk00000001_sig00000543,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1b
    );
  blk00000001_blk000005a6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000542,
      I1 => blk00000001_sig00000543,
      I2 => blk00000001_sig00000543,
      I3 => blk00000001_sig00000543,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a1a
    );
  blk00000001_blk000005a5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000541,
      I1 => blk00000001_sig00000542,
      I2 => blk00000001_sig00000543,
      I3 => blk00000001_sig00000543,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a19
    );
  blk00000001_blk000005a4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000540,
      I1 => blk00000001_sig00000541,
      I2 => blk00000001_sig00000542,
      I3 => blk00000001_sig00000543,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a18
    );
  blk00000001_blk000005a3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053f,
      I1 => blk00000001_sig00000540,
      I2 => blk00000001_sig00000541,
      I3 => blk00000001_sig00000542,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a17
    );
  blk00000001_blk000005a2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053e,
      I1 => blk00000001_sig0000053f,
      I2 => blk00000001_sig00000540,
      I3 => blk00000001_sig00000541,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a16
    );
  blk00000001_blk000005a1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053d,
      I1 => blk00000001_sig0000053e,
      I2 => blk00000001_sig0000053f,
      I3 => blk00000001_sig00000540,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a15
    );
  blk00000001_blk000005a0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053c,
      I1 => blk00000001_sig0000053d,
      I2 => blk00000001_sig0000053e,
      I3 => blk00000001_sig0000053f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a14
    );
  blk00000001_blk0000059f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053b,
      I1 => blk00000001_sig0000053c,
      I2 => blk00000001_sig0000053d,
      I3 => blk00000001_sig0000053e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a13
    );
  blk00000001_blk0000059e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000053a,
      I1 => blk00000001_sig0000053b,
      I2 => blk00000001_sig0000053c,
      I3 => blk00000001_sig0000053d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a12
    );
  blk00000001_blk0000059d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000539,
      I1 => blk00000001_sig0000053a,
      I2 => blk00000001_sig0000053b,
      I3 => blk00000001_sig0000053c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a11
    );
  blk00000001_blk0000059c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000538,
      I1 => blk00000001_sig00000539,
      I2 => blk00000001_sig0000053a,
      I3 => blk00000001_sig0000053b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a10
    );
  blk00000001_blk0000059b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000537,
      I1 => blk00000001_sig00000538,
      I2 => blk00000001_sig00000539,
      I3 => blk00000001_sig0000053a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0f
    );
  blk00000001_blk0000059a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000536,
      I1 => blk00000001_sig00000537,
      I2 => blk00000001_sig00000538,
      I3 => blk00000001_sig00000539,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0e
    );
  blk00000001_blk00000599 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000535,
      I1 => blk00000001_sig00000536,
      I2 => blk00000001_sig00000537,
      I3 => blk00000001_sig00000538,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0d
    );
  blk00000001_blk00000598 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000534,
      I1 => blk00000001_sig00000535,
      I2 => blk00000001_sig00000536,
      I3 => blk00000001_sig00000537,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0c
    );
  blk00000001_blk00000597 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000533,
      I1 => blk00000001_sig00000534,
      I2 => blk00000001_sig00000535,
      I3 => blk00000001_sig00000536,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0b
    );
  blk00000001_blk00000596 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000532,
      I1 => blk00000001_sig00000533,
      I2 => blk00000001_sig00000534,
      I3 => blk00000001_sig00000535,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a0a
    );
  blk00000001_blk00000595 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000531,
      I1 => blk00000001_sig00000532,
      I2 => blk00000001_sig00000533,
      I3 => blk00000001_sig00000534,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a09
    );
  blk00000001_blk00000594 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000530,
      I1 => blk00000001_sig00000531,
      I2 => blk00000001_sig00000532,
      I3 => blk00000001_sig00000533,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a08
    );
  blk00000001_blk00000593 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052f,
      I1 => blk00000001_sig00000530,
      I2 => blk00000001_sig00000531,
      I3 => blk00000001_sig00000532,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a07
    );
  blk00000001_blk00000592 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000052e,
      I1 => blk00000001_sig0000052f,
      I2 => blk00000001_sig00000530,
      I3 => blk00000001_sig00000531,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a06
    );
  blk00000001_blk00000591 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig0000052e,
      I2 => blk00000001_sig0000052f,
      I3 => blk00000001_sig00000530,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a05
    );
  blk00000001_blk00000590 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig0000052e,
      I3 => blk00000001_sig0000052f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a04
    );
  blk00000001_blk0000058f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig0000052e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a03
    );
  blk00000001_blk0000058e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a02,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d1
    );
  blk00000001_blk0000058d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a01,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d0
    );
  blk00000001_blk0000058c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000a00,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006cf
    );
  blk00000001_blk0000058b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ff,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a7
    );
  blk00000001_blk0000058a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009fe,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a6
    );
  blk00000001_blk00000589 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009fd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a5
    );
  blk00000001_blk00000588 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009fc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a4
    );
  blk00000001_blk00000587 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009fb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a3
    );
  blk00000001_blk00000586 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009fa,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a2
    );
  blk00000001_blk00000585 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a1
    );
  blk00000001_blk00000584 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a0
    );
  blk00000001_blk00000583 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039f
    );
  blk00000001_blk00000582 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039e
    );
  blk00000001_blk00000581 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039d
    );
  blk00000001_blk00000580 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039c
    );
  blk00000001_blk0000057f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039b
    );
  blk00000001_blk0000057e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000039a
    );
  blk00000001_blk0000057d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000399
    );
  blk00000001_blk0000057c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009f0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000398
    );
  blk00000001_blk0000057b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ef,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000057b_Q_UNCONNECTED
    );
  blk00000001_blk0000057a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ee,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk0000057a_Q_UNCONNECTED
    );
  blk00000001_blk00000579 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ed,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000579_Q_UNCONNECTED
    );
  blk00000001_blk00000578 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ec,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000578_Q_UNCONNECTED
    );
  blk00000001_blk00000577 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009eb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000577_Q_UNCONNECTED
    );
  blk00000001_blk00000576 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ea,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000576_Q_UNCONNECTED
    );
  blk00000001_blk00000575 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000559,
      I1 => blk00000001_sig00000559,
      I2 => blk00000001_sig00000559,
      I3 => blk00000001_sig00000559,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a02
    );
  blk00000001_blk00000574 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000558,
      I1 => blk00000001_sig00000559,
      I2 => blk00000001_sig00000559,
      I3 => blk00000001_sig00000559,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a01
    );
  blk00000001_blk00000573 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000557,
      I1 => blk00000001_sig00000558,
      I2 => blk00000001_sig00000559,
      I3 => blk00000001_sig00000559,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000a00
    );
  blk00000001_blk00000572 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000556,
      I1 => blk00000001_sig00000557,
      I2 => blk00000001_sig00000558,
      I3 => blk00000001_sig00000559,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ff
    );
  blk00000001_blk00000571 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000555,
      I1 => blk00000001_sig00000556,
      I2 => blk00000001_sig00000557,
      I3 => blk00000001_sig00000558,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009fe
    );
  blk00000001_blk00000570 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000554,
      I1 => blk00000001_sig00000555,
      I2 => blk00000001_sig00000556,
      I3 => blk00000001_sig00000557,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009fd
    );
  blk00000001_blk0000056f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000553,
      I1 => blk00000001_sig00000554,
      I2 => blk00000001_sig00000555,
      I3 => blk00000001_sig00000556,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009fc
    );
  blk00000001_blk0000056e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000552,
      I1 => blk00000001_sig00000553,
      I2 => blk00000001_sig00000554,
      I3 => blk00000001_sig00000555,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009fb
    );
  blk00000001_blk0000056d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000551,
      I1 => blk00000001_sig00000552,
      I2 => blk00000001_sig00000553,
      I3 => blk00000001_sig00000554,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009fa
    );
  blk00000001_blk0000056c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000550,
      I1 => blk00000001_sig00000551,
      I2 => blk00000001_sig00000552,
      I3 => blk00000001_sig00000553,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f9
    );
  blk00000001_blk0000056b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054f,
      I1 => blk00000001_sig00000550,
      I2 => blk00000001_sig00000551,
      I3 => blk00000001_sig00000552,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f8
    );
  blk00000001_blk0000056a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054e,
      I1 => blk00000001_sig0000054f,
      I2 => blk00000001_sig00000550,
      I3 => blk00000001_sig00000551,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f7
    );
  blk00000001_blk00000569 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054d,
      I1 => blk00000001_sig0000054e,
      I2 => blk00000001_sig0000054f,
      I3 => blk00000001_sig00000550,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f6
    );
  blk00000001_blk00000568 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054c,
      I1 => blk00000001_sig0000054d,
      I2 => blk00000001_sig0000054e,
      I3 => blk00000001_sig0000054f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f5
    );
  blk00000001_blk00000567 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054b,
      I1 => blk00000001_sig0000054c,
      I2 => blk00000001_sig0000054d,
      I3 => blk00000001_sig0000054e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f4
    );
  blk00000001_blk00000566 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000054a,
      I1 => blk00000001_sig0000054b,
      I2 => blk00000001_sig0000054c,
      I3 => blk00000001_sig0000054d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f3
    );
  blk00000001_blk00000565 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000549,
      I1 => blk00000001_sig0000054a,
      I2 => blk00000001_sig0000054b,
      I3 => blk00000001_sig0000054c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f2
    );
  blk00000001_blk00000564 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000548,
      I1 => blk00000001_sig00000549,
      I2 => blk00000001_sig0000054a,
      I3 => blk00000001_sig0000054b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f1
    );
  blk00000001_blk00000563 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000547,
      I1 => blk00000001_sig00000548,
      I2 => blk00000001_sig00000549,
      I3 => blk00000001_sig0000054a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009f0
    );
  blk00000001_blk00000562 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000546,
      I1 => blk00000001_sig00000547,
      I2 => blk00000001_sig00000548,
      I3 => blk00000001_sig00000549,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ef
    );
  blk00000001_blk00000561 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000545,
      I1 => blk00000001_sig00000546,
      I2 => blk00000001_sig00000547,
      I3 => blk00000001_sig00000548,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ee
    );
  blk00000001_blk00000560 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000544,
      I1 => blk00000001_sig00000545,
      I2 => blk00000001_sig00000546,
      I3 => blk00000001_sig00000547,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ed
    );
  blk00000001_blk0000055f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000544,
      I2 => blk00000001_sig00000545,
      I3 => blk00000001_sig00000546,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ec
    );
  blk00000001_blk0000055e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000544,
      I3 => blk00000001_sig00000545,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009eb
    );
  blk00000001_blk0000055d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig00000544,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ea
    );
  blk00000001_blk0000055c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d4
    );
  blk00000001_blk0000055b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d3
    );
  blk00000001_blk0000055a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d2
    );
  blk00000001_blk00000559 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b7
    );
  blk00000001_blk00000558 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b6
    );
  blk00000001_blk00000557 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b5
    );
  blk00000001_blk00000556 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b4
    );
  blk00000001_blk00000555 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b3
    );
  blk00000001_blk00000554 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b2
    );
  blk00000001_blk00000553 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009e0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b1
    );
  blk00000001_blk00000552 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009df,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b0
    );
  blk00000001_blk00000551 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009de,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003af
    );
  blk00000001_blk00000550 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009dd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ae
    );
  blk00000001_blk0000054f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009dc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ad
    );
  blk00000001_blk0000054e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009db,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ac
    );
  blk00000001_blk0000054d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009da,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ab
    );
  blk00000001_blk0000054c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003aa
    );
  blk00000001_blk0000054b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a9
    );
  blk00000001_blk0000054a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003a8
    );
  blk00000001_blk00000549 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000549_Q_UNCONNECTED
    );
  blk00000001_blk00000548 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000548_Q_UNCONNECTED
    );
  blk00000001_blk00000547 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000547_Q_UNCONNECTED
    );
  blk00000001_blk00000546 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000546_Q_UNCONNECTED
    );
  blk00000001_blk00000545 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000545_Q_UNCONNECTED
    );
  blk00000001_blk00000544 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000544_Q_UNCONNECTED
    );
  blk00000001_blk00000543 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056f,
      I1 => blk00000001_sig0000056f,
      I2 => blk00000001_sig0000056f,
      I3 => blk00000001_sig0000056f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e9
    );
  blk00000001_blk00000542 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056e,
      I1 => blk00000001_sig0000056f,
      I2 => blk00000001_sig0000056f,
      I3 => blk00000001_sig0000056f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e8
    );
  blk00000001_blk00000541 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056d,
      I1 => blk00000001_sig0000056e,
      I2 => blk00000001_sig0000056f,
      I3 => blk00000001_sig0000056f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e7
    );
  blk00000001_blk00000540 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056c,
      I1 => blk00000001_sig0000056d,
      I2 => blk00000001_sig0000056e,
      I3 => blk00000001_sig0000056f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e6
    );
  blk00000001_blk0000053f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056b,
      I1 => blk00000001_sig0000056c,
      I2 => blk00000001_sig0000056d,
      I3 => blk00000001_sig0000056e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e5
    );
  blk00000001_blk0000053e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000056a,
      I1 => blk00000001_sig0000056b,
      I2 => blk00000001_sig0000056c,
      I3 => blk00000001_sig0000056d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e4
    );
  blk00000001_blk0000053d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000569,
      I1 => blk00000001_sig0000056a,
      I2 => blk00000001_sig0000056b,
      I3 => blk00000001_sig0000056c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e3
    );
  blk00000001_blk0000053c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000568,
      I1 => blk00000001_sig00000569,
      I2 => blk00000001_sig0000056a,
      I3 => blk00000001_sig0000056b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e2
    );
  blk00000001_blk0000053b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000567,
      I1 => blk00000001_sig00000568,
      I2 => blk00000001_sig00000569,
      I3 => blk00000001_sig0000056a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e1
    );
  blk00000001_blk0000053a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000566,
      I1 => blk00000001_sig00000567,
      I2 => blk00000001_sig00000568,
      I3 => blk00000001_sig00000569,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009e0
    );
  blk00000001_blk00000539 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000565,
      I1 => blk00000001_sig00000566,
      I2 => blk00000001_sig00000567,
      I3 => blk00000001_sig00000568,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009df
    );
  blk00000001_blk00000538 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000564,
      I1 => blk00000001_sig00000565,
      I2 => blk00000001_sig00000566,
      I3 => blk00000001_sig00000567,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009de
    );
  blk00000001_blk00000537 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000563,
      I1 => blk00000001_sig00000564,
      I2 => blk00000001_sig00000565,
      I3 => blk00000001_sig00000566,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009dd
    );
  blk00000001_blk00000536 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000562,
      I1 => blk00000001_sig00000563,
      I2 => blk00000001_sig00000564,
      I3 => blk00000001_sig00000565,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009dc
    );
  blk00000001_blk00000535 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000561,
      I1 => blk00000001_sig00000562,
      I2 => blk00000001_sig00000563,
      I3 => blk00000001_sig00000564,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009db
    );
  blk00000001_blk00000534 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000560,
      I1 => blk00000001_sig00000561,
      I2 => blk00000001_sig00000562,
      I3 => blk00000001_sig00000563,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009da
    );
  blk00000001_blk00000533 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055f,
      I1 => blk00000001_sig00000560,
      I2 => blk00000001_sig00000561,
      I3 => blk00000001_sig00000562,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d9
    );
  blk00000001_blk00000532 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055e,
      I1 => blk00000001_sig0000055f,
      I2 => blk00000001_sig00000560,
      I3 => blk00000001_sig00000561,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d8
    );
  blk00000001_blk00000531 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055d,
      I1 => blk00000001_sig0000055e,
      I2 => blk00000001_sig0000055f,
      I3 => blk00000001_sig00000560,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d7
    );
  blk00000001_blk00000530 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055c,
      I1 => blk00000001_sig0000055d,
      I2 => blk00000001_sig0000055e,
      I3 => blk00000001_sig0000055f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d6
    );
  blk00000001_blk0000052f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055b,
      I1 => blk00000001_sig0000055c,
      I2 => blk00000001_sig0000055d,
      I3 => blk00000001_sig0000055e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d5
    );
  blk00000001_blk0000052e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000055a,
      I1 => blk00000001_sig0000055b,
      I2 => blk00000001_sig0000055c,
      I3 => blk00000001_sig0000055d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d4
    );
  blk00000001_blk0000052d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig0000055a,
      I2 => blk00000001_sig0000055b,
      I3 => blk00000001_sig0000055c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d3
    );
  blk00000001_blk0000052c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig0000055a,
      I3 => blk00000001_sig0000055b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d2
    );
  blk00000001_blk0000052b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig0000055a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d1
    );
  blk00000001_blk0000052a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009d0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d7
    );
  blk00000001_blk00000529 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009cf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d6
    );
  blk00000001_blk00000528 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ce,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d5
    );
  blk00000001_blk00000527 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009cd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c7
    );
  blk00000001_blk00000526 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009cc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c6
    );
  blk00000001_blk00000525 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009cb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c5
    );
  blk00000001_blk00000524 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ca,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c4
    );
  blk00000001_blk00000523 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c3
    );
  blk00000001_blk00000522 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c2
    );
  blk00000001_blk00000521 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c1
    );
  blk00000001_blk00000520 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c0
    );
  blk00000001_blk0000051f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003bf
    );
  blk00000001_blk0000051e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003be
    );
  blk00000001_blk0000051d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003bd
    );
  blk00000001_blk0000051c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003bc
    );
  blk00000001_blk0000051b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003bb
    );
  blk00000001_blk0000051a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009c0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ba
    );
  blk00000001_blk00000519 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009bf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b9
    );
  blk00000001_blk00000518 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009be,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003b8
    );
  blk00000001_blk00000517 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009bd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000517_Q_UNCONNECTED
    );
  blk00000001_blk00000516 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009bc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000516_Q_UNCONNECTED
    );
  blk00000001_blk00000515 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009bb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000515_Q_UNCONNECTED
    );
  blk00000001_blk00000514 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ba,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000514_Q_UNCONNECTED
    );
  blk00000001_blk00000513 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000513_Q_UNCONNECTED
    );
  blk00000001_blk00000512 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk00000512_Q_UNCONNECTED
    );
  blk00000001_blk00000511 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000585,
      I1 => blk00000001_sig00000585,
      I2 => blk00000001_sig00000585,
      I3 => blk00000001_sig00000585,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009d0
    );
  blk00000001_blk00000510 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000584,
      I1 => blk00000001_sig00000585,
      I2 => blk00000001_sig00000585,
      I3 => blk00000001_sig00000585,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009cf
    );
  blk00000001_blk0000050f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000583,
      I1 => blk00000001_sig00000584,
      I2 => blk00000001_sig00000585,
      I3 => blk00000001_sig00000585,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ce
    );
  blk00000001_blk0000050e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000582,
      I1 => blk00000001_sig00000583,
      I2 => blk00000001_sig00000584,
      I3 => blk00000001_sig00000585,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009cd
    );
  blk00000001_blk0000050d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000581,
      I1 => blk00000001_sig00000582,
      I2 => blk00000001_sig00000583,
      I3 => blk00000001_sig00000584,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009cc
    );
  blk00000001_blk0000050c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000580,
      I1 => blk00000001_sig00000581,
      I2 => blk00000001_sig00000582,
      I3 => blk00000001_sig00000583,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009cb
    );
  blk00000001_blk0000050b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057f,
      I1 => blk00000001_sig00000580,
      I2 => blk00000001_sig00000581,
      I3 => blk00000001_sig00000582,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ca
    );
  blk00000001_blk0000050a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057e,
      I1 => blk00000001_sig0000057f,
      I2 => blk00000001_sig00000580,
      I3 => blk00000001_sig00000581,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c9
    );
  blk00000001_blk00000509 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057d,
      I1 => blk00000001_sig0000057e,
      I2 => blk00000001_sig0000057f,
      I3 => blk00000001_sig00000580,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c8
    );
  blk00000001_blk00000508 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057c,
      I1 => blk00000001_sig0000057d,
      I2 => blk00000001_sig0000057e,
      I3 => blk00000001_sig0000057f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c7
    );
  blk00000001_blk00000507 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057b,
      I1 => blk00000001_sig0000057c,
      I2 => blk00000001_sig0000057d,
      I3 => blk00000001_sig0000057e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c6
    );
  blk00000001_blk00000506 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000057a,
      I1 => blk00000001_sig0000057b,
      I2 => blk00000001_sig0000057c,
      I3 => blk00000001_sig0000057d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c5
    );
  blk00000001_blk00000505 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000579,
      I1 => blk00000001_sig0000057a,
      I2 => blk00000001_sig0000057b,
      I3 => blk00000001_sig0000057c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c4
    );
  blk00000001_blk00000504 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000578,
      I1 => blk00000001_sig00000579,
      I2 => blk00000001_sig0000057a,
      I3 => blk00000001_sig0000057b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c3
    );
  blk00000001_blk00000503 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000577,
      I1 => blk00000001_sig00000578,
      I2 => blk00000001_sig00000579,
      I3 => blk00000001_sig0000057a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c2
    );
  blk00000001_blk00000502 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000576,
      I1 => blk00000001_sig00000577,
      I2 => blk00000001_sig00000578,
      I3 => blk00000001_sig00000579,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c1
    );
  blk00000001_blk00000501 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000575,
      I1 => blk00000001_sig00000576,
      I2 => blk00000001_sig00000577,
      I3 => blk00000001_sig00000578,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009c0
    );
  blk00000001_blk00000500 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000574,
      I1 => blk00000001_sig00000575,
      I2 => blk00000001_sig00000576,
      I3 => blk00000001_sig00000577,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009bf
    );
  blk00000001_blk000004ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000573,
      I1 => blk00000001_sig00000574,
      I2 => blk00000001_sig00000575,
      I3 => blk00000001_sig00000576,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009be
    );
  blk00000001_blk000004fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000572,
      I1 => blk00000001_sig00000573,
      I2 => blk00000001_sig00000574,
      I3 => blk00000001_sig00000575,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009bd
    );
  blk00000001_blk000004fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000571,
      I1 => blk00000001_sig00000572,
      I2 => blk00000001_sig00000573,
      I3 => blk00000001_sig00000574,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009bc
    );
  blk00000001_blk000004fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000570,
      I1 => blk00000001_sig00000571,
      I2 => blk00000001_sig00000572,
      I3 => blk00000001_sig00000573,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009bb
    );
  blk00000001_blk000004fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000570,
      I2 => blk00000001_sig00000571,
      I3 => blk00000001_sig00000572,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ba
    );
  blk00000001_blk000004fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000570,
      I3 => blk00000001_sig00000571,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b9
    );
  blk00000001_blk000004f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig00000570,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b8
    );
  blk00000001_blk000004f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006da
    );
  blk00000001_blk000004f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d9
    );
  blk00000001_blk000004f6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006d8
    );
  blk00000001_blk000004f5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d7
    );
  blk00000001_blk000004f4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d6
    );
  blk00000001_blk000004f3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d5
    );
  blk00000001_blk000004f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d4
    );
  blk00000001_blk000004f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009b0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d3
    );
  blk00000001_blk000004f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009af,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d2
    );
  blk00000001_blk000004ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ae,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d1
    );
  blk00000001_blk000004ee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ad,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d0
    );
  blk00000001_blk000004ed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ac,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003cf
    );
  blk00000001_blk000004ec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009ab,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ce
    );
  blk00000001_blk000004eb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009aa,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003cd
    );
  blk00000001_blk000004ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003cc
    );
  blk00000001_blk000004e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003cb
    );
  blk00000001_blk000004e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003ca
    );
  blk00000001_blk000004e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c9
    );
  blk00000001_blk000004e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003c8
    );
  blk00000001_blk000004e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e5_Q_UNCONNECTED
    );
  blk00000001_blk000004e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e4_Q_UNCONNECTED
    );
  blk00000001_blk000004e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e3_Q_UNCONNECTED
    );
  blk00000001_blk000004e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e2_Q_UNCONNECTED
    );
  blk00000001_blk000004e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000009a0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e1_Q_UNCONNECTED
    );
  blk00000001_blk000004e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004e0_Q_UNCONNECTED
    );
  blk00000001_blk000004df : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059b,
      I1 => blk00000001_sig0000059b,
      I2 => blk00000001_sig0000059b,
      I3 => blk00000001_sig0000059b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b7
    );
  blk00000001_blk000004de : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059a,
      I1 => blk00000001_sig0000059b,
      I2 => blk00000001_sig0000059b,
      I3 => blk00000001_sig0000059b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b6
    );
  blk00000001_blk000004dd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000599,
      I1 => blk00000001_sig0000059a,
      I2 => blk00000001_sig0000059b,
      I3 => blk00000001_sig0000059b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b5
    );
  blk00000001_blk000004dc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000598,
      I1 => blk00000001_sig00000599,
      I2 => blk00000001_sig0000059a,
      I3 => blk00000001_sig0000059b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b4
    );
  blk00000001_blk000004db : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000597,
      I1 => blk00000001_sig00000598,
      I2 => blk00000001_sig00000599,
      I3 => blk00000001_sig0000059a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b3
    );
  blk00000001_blk000004da : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000596,
      I1 => blk00000001_sig00000597,
      I2 => blk00000001_sig00000598,
      I3 => blk00000001_sig00000599,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b2
    );
  blk00000001_blk000004d9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000595,
      I1 => blk00000001_sig00000596,
      I2 => blk00000001_sig00000597,
      I3 => blk00000001_sig00000598,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b1
    );
  blk00000001_blk000004d8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000594,
      I1 => blk00000001_sig00000595,
      I2 => blk00000001_sig00000596,
      I3 => blk00000001_sig00000597,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009b0
    );
  blk00000001_blk000004d7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000593,
      I1 => blk00000001_sig00000594,
      I2 => blk00000001_sig00000595,
      I3 => blk00000001_sig00000596,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009af
    );
  blk00000001_blk000004d6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000592,
      I1 => blk00000001_sig00000593,
      I2 => blk00000001_sig00000594,
      I3 => blk00000001_sig00000595,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ae
    );
  blk00000001_blk000004d5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000591,
      I1 => blk00000001_sig00000592,
      I2 => blk00000001_sig00000593,
      I3 => blk00000001_sig00000594,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ad
    );
  blk00000001_blk000004d4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000590,
      I1 => blk00000001_sig00000591,
      I2 => blk00000001_sig00000592,
      I3 => blk00000001_sig00000593,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ac
    );
  blk00000001_blk000004d3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058f,
      I1 => blk00000001_sig00000590,
      I2 => blk00000001_sig00000591,
      I3 => blk00000001_sig00000592,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009ab
    );
  blk00000001_blk000004d2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058e,
      I1 => blk00000001_sig0000058f,
      I2 => blk00000001_sig00000590,
      I3 => blk00000001_sig00000591,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009aa
    );
  blk00000001_blk000004d1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058d,
      I1 => blk00000001_sig0000058e,
      I2 => blk00000001_sig0000058f,
      I3 => blk00000001_sig00000590,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a9
    );
  blk00000001_blk000004d0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058c,
      I1 => blk00000001_sig0000058d,
      I2 => blk00000001_sig0000058e,
      I3 => blk00000001_sig0000058f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a8
    );
  blk00000001_blk000004cf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058b,
      I1 => blk00000001_sig0000058c,
      I2 => blk00000001_sig0000058d,
      I3 => blk00000001_sig0000058e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a7
    );
  blk00000001_blk000004ce : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000058a,
      I1 => blk00000001_sig0000058b,
      I2 => blk00000001_sig0000058c,
      I3 => blk00000001_sig0000058d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a6
    );
  blk00000001_blk000004cd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000589,
      I1 => blk00000001_sig0000058a,
      I2 => blk00000001_sig0000058b,
      I3 => blk00000001_sig0000058c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a5
    );
  blk00000001_blk000004cc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000588,
      I1 => blk00000001_sig00000589,
      I2 => blk00000001_sig0000058a,
      I3 => blk00000001_sig0000058b,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a4
    );
  blk00000001_blk000004cb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000587,
      I1 => blk00000001_sig00000588,
      I2 => blk00000001_sig00000589,
      I3 => blk00000001_sig0000058a,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a3
    );
  blk00000001_blk000004ca : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000586,
      I1 => blk00000001_sig00000587,
      I2 => blk00000001_sig00000588,
      I3 => blk00000001_sig00000589,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a2
    );
  blk00000001_blk000004c9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig00000586,
      I2 => blk00000001_sig00000587,
      I3 => blk00000001_sig00000588,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a1
    );
  blk00000001_blk000004c8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig00000586,
      I3 => blk00000001_sig00000587,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig000009a0
    );
  blk00000001_blk000004c7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig00000586,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099f
    );
  blk00000001_blk000004c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006dd
    );
  blk00000001_blk000004c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006dc
    );
  blk00000001_blk000004c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000006db
    );
  blk00000001_blk000004c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e7
    );
  blk00000001_blk000004c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000099a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e6
    );
  blk00000001_blk000004c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000999,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e5
    );
  blk00000001_blk000004c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000998,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e4
    );
  blk00000001_blk000004bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000997,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e3
    );
  blk00000001_blk000004be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000996,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e2
    );
  blk00000001_blk000004bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000995,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e1
    );
  blk00000001_blk000004bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000994,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003e0
    );
  blk00000001_blk000004bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000993,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003df
    );
  blk00000001_blk000004ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000992,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003de
    );
  blk00000001_blk000004b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000991,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003dd
    );
  blk00000001_blk000004b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000990,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003dc
    );
  blk00000001_blk000004b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003db
    );
  blk00000001_blk000004b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003da
    );
  blk00000001_blk000004b5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d9
    );
  blk00000001_blk000004b4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000003d8
    );
  blk00000001_blk000004b3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004b3_Q_UNCONNECTED
    );
  blk00000001_blk000004b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000098a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004b2_Q_UNCONNECTED
    );
  blk00000001_blk000004b1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000989,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004b1_Q_UNCONNECTED
    );
  blk00000001_blk000004b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000988,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004b0_Q_UNCONNECTED
    );
  blk00000001_blk000004af : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000987,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004af_Q_UNCONNECTED
    );
  blk00000001_blk000004ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000986,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => NLW_blk00000001_blk000004ae_Q_UNCONNECTED
    );
  blk00000001_blk000004ad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005b1,
      I1 => blk00000001_sig000005b1,
      I2 => blk00000001_sig000005b1,
      I3 => blk00000001_sig000005b1,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099e
    );
  blk00000001_blk000004ac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005b0,
      I1 => blk00000001_sig000005b1,
      I2 => blk00000001_sig000005b1,
      I3 => blk00000001_sig000005b1,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099d
    );
  blk00000001_blk000004ab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005af,
      I1 => blk00000001_sig000005b0,
      I2 => blk00000001_sig000005b1,
      I3 => blk00000001_sig000005b1,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099c
    );
  blk00000001_blk000004aa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005ae,
      I1 => blk00000001_sig000005af,
      I2 => blk00000001_sig000005b0,
      I3 => blk00000001_sig000005b1,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099b
    );
  blk00000001_blk000004a9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005ad,
      I1 => blk00000001_sig000005ae,
      I2 => blk00000001_sig000005af,
      I3 => blk00000001_sig000005b0,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000099a
    );
  blk00000001_blk000004a8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005ac,
      I1 => blk00000001_sig000005ad,
      I2 => blk00000001_sig000005ae,
      I3 => blk00000001_sig000005af,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000999
    );
  blk00000001_blk000004a7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005ab,
      I1 => blk00000001_sig000005ac,
      I2 => blk00000001_sig000005ad,
      I3 => blk00000001_sig000005ae,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000998
    );
  blk00000001_blk000004a6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005aa,
      I1 => blk00000001_sig000005ab,
      I2 => blk00000001_sig000005ac,
      I3 => blk00000001_sig000005ad,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000997
    );
  blk00000001_blk000004a5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a9,
      I1 => blk00000001_sig000005aa,
      I2 => blk00000001_sig000005ab,
      I3 => blk00000001_sig000005ac,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000996
    );
  blk00000001_blk000004a4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a8,
      I1 => blk00000001_sig000005a9,
      I2 => blk00000001_sig000005aa,
      I3 => blk00000001_sig000005ab,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000995
    );
  blk00000001_blk000004a3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a7,
      I1 => blk00000001_sig000005a8,
      I2 => blk00000001_sig000005a9,
      I3 => blk00000001_sig000005aa,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000994
    );
  blk00000001_blk000004a2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a6,
      I1 => blk00000001_sig000005a7,
      I2 => blk00000001_sig000005a8,
      I3 => blk00000001_sig000005a9,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000993
    );
  blk00000001_blk000004a1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a5,
      I1 => blk00000001_sig000005a6,
      I2 => blk00000001_sig000005a7,
      I3 => blk00000001_sig000005a8,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000992
    );
  blk00000001_blk000004a0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a4,
      I1 => blk00000001_sig000005a5,
      I2 => blk00000001_sig000005a6,
      I3 => blk00000001_sig000005a7,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000991
    );
  blk00000001_blk0000049f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a3,
      I1 => blk00000001_sig000005a4,
      I2 => blk00000001_sig000005a5,
      I3 => blk00000001_sig000005a6,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000990
    );
  blk00000001_blk0000049e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a2,
      I1 => blk00000001_sig000005a3,
      I2 => blk00000001_sig000005a4,
      I3 => blk00000001_sig000005a5,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098f
    );
  blk00000001_blk0000049d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a1,
      I1 => blk00000001_sig000005a2,
      I2 => blk00000001_sig000005a3,
      I3 => blk00000001_sig000005a4,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098e
    );
  blk00000001_blk0000049c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000005a0,
      I1 => blk00000001_sig000005a1,
      I2 => blk00000001_sig000005a2,
      I3 => blk00000001_sig000005a3,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098d
    );
  blk00000001_blk0000049b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059f,
      I1 => blk00000001_sig000005a0,
      I2 => blk00000001_sig000005a1,
      I3 => blk00000001_sig000005a2,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098c
    );
  blk00000001_blk0000049a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059e,
      I1 => blk00000001_sig0000059f,
      I2 => blk00000001_sig000005a0,
      I3 => blk00000001_sig000005a1,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098b
    );
  blk00000001_blk00000499 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059d,
      I1 => blk00000001_sig0000059e,
      I2 => blk00000001_sig0000059f,
      I3 => blk00000001_sig000005a0,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig0000098a
    );
  blk00000001_blk00000498 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000059c,
      I1 => blk00000001_sig0000059d,
      I2 => blk00000001_sig0000059e,
      I3 => blk00000001_sig0000059f,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000989
    );
  blk00000001_blk00000497 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => blk00000001_sig0000059c,
      I2 => blk00000001_sig0000059d,
      I3 => blk00000001_sig0000059e,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000988
    );
  blk00000001_blk00000496 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => blk00000001_sig0000059c,
      I3 => blk00000001_sig0000059d,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000987
    );
  blk00000001_blk00000495 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      I3 => blk00000001_sig0000059c,
      I4 => blk00000001_sig000002e5,
      I5 => blk00000001_sig000002e6,
      O => blk00000001_sig00000986
    );
  blk00000001_blk00000494 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000008af,
      Q => blk00000001_sig00000985
    );
  blk00000001_blk00000493 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001e0,
      Q => blk00000001_sig00000922
    );
  blk00000001_blk00000492 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000922,
      Q => blk00000001_sig000007c7
    );
  blk00000001_blk00000491 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000da6,
      Q => blk00000001_sig000008af
    );
  blk00000001_blk00000490 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000001d9,
      Q => blk00000001_sig00000984
    );
  blk00000001_blk0000048f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000984,
      Q => blk00000001_sig000008ae
    );
  blk00000001_blk0000048e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000795,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000766
    );
  blk00000001_blk0000048d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000794,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000767
    );
  blk00000001_blk0000048c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000793,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000768
    );
  blk00000001_blk0000048b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000792,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000769
    );
  blk00000001_blk0000048a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000791,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076a
    );
  blk00000001_blk00000489 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000790,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076b
    );
  blk00000001_blk00000488 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076c
    );
  blk00000001_blk00000487 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076d
    );
  blk00000001_blk00000486 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076e
    );
  blk00000001_blk00000485 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000076f
    );
  blk00000001_blk00000484 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000770
    );
  blk00000001_blk00000483 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000078a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000771
    );
  blk00000001_blk00000482 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000789,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000772
    );
  blk00000001_blk00000481 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000788,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000773
    );
  blk00000001_blk00000480 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000787,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000774
    );
  blk00000001_blk0000047f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000786,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000775
    );
  blk00000001_blk0000047e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f8,
      Q => blk00000001_sig00000795
    );
  blk00000001_blk0000047d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f9,
      Q => blk00000001_sig00000794
    );
  blk00000001_blk0000047c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003fa,
      Q => blk00000001_sig00000793
    );
  blk00000001_blk0000047b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003fb,
      Q => blk00000001_sig00000792
    );
  blk00000001_blk0000047a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003fc,
      Q => blk00000001_sig00000791
    );
  blk00000001_blk00000479 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003fd,
      Q => blk00000001_sig00000790
    );
  blk00000001_blk00000478 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003fe,
      Q => blk00000001_sig0000078f
    );
  blk00000001_blk00000477 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ff,
      Q => blk00000001_sig0000078e
    );
  blk00000001_blk00000476 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000400,
      Q => blk00000001_sig0000078d
    );
  blk00000001_blk00000475 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000401,
      Q => blk00000001_sig0000078c
    );
  blk00000001_blk00000474 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000402,
      Q => blk00000001_sig0000078b
    );
  blk00000001_blk00000473 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000403,
      Q => blk00000001_sig0000078a
    );
  blk00000001_blk00000472 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000404,
      Q => blk00000001_sig00000789
    );
  blk00000001_blk00000471 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000405,
      Q => blk00000001_sig00000788
    );
  blk00000001_blk00000470 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000406,
      Q => blk00000001_sig00000787
    );
  blk00000001_blk0000046f : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000407,
      Q => blk00000001_sig00000786
    );
  blk00000001_blk0000046e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000785,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000756
    );
  blk00000001_blk0000046d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000784,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000757
    );
  blk00000001_blk0000046c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000783,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000758
    );
  blk00000001_blk0000046b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000782,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000759
    );
  blk00000001_blk0000046a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000781,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075a
    );
  blk00000001_blk00000469 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000780,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075b
    );
  blk00000001_blk00000468 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075c
    );
  blk00000001_blk00000467 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075d
    );
  blk00000001_blk00000466 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075e
    );
  blk00000001_blk00000465 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000075f
    );
  blk00000001_blk00000464 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000760
    );
  blk00000001_blk00000463 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000077a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000761
    );
  blk00000001_blk00000462 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000779,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000762
    );
  blk00000001_blk00000461 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000778,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000763
    );
  blk00000001_blk00000460 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000777,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000764
    );
  blk00000001_blk0000045f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000776,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000765
    );
  blk00000001_blk0000045e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003e8,
      Q => blk00000001_sig00000785
    );
  blk00000001_blk0000045d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003e9,
      Q => blk00000001_sig00000784
    );
  blk00000001_blk0000045c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ea,
      Q => blk00000001_sig00000783
    );
  blk00000001_blk0000045b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003eb,
      Q => blk00000001_sig00000782
    );
  blk00000001_blk0000045a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ec,
      Q => blk00000001_sig00000781
    );
  blk00000001_blk00000459 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ed,
      Q => blk00000001_sig00000780
    );
  blk00000001_blk00000458 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ee,
      Q => blk00000001_sig0000077f
    );
  blk00000001_blk00000457 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003ef,
      Q => blk00000001_sig0000077e
    );
  blk00000001_blk00000456 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f0,
      Q => blk00000001_sig0000077d
    );
  blk00000001_blk00000455 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f1,
      Q => blk00000001_sig0000077c
    );
  blk00000001_blk00000454 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f2,
      Q => blk00000001_sig0000077b
    );
  blk00000001_blk00000453 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f3,
      Q => blk00000001_sig0000077a
    );
  blk00000001_blk00000452 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f4,
      Q => blk00000001_sig00000779
    );
  blk00000001_blk00000451 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f5,
      Q => blk00000001_sig00000778
    );
  blk00000001_blk00000450 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f6,
      Q => blk00000001_sig00000777
    );
  blk00000001_blk0000044f : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => blk00000001_sig000000c0,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000003f7,
      Q => blk00000001_sig00000776
    );
  blk00000001_blk0000044e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072e,
      Q => blk00000001_sig00000602
    );
  blk00000001_blk0000044d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072f,
      Q => blk00000001_sig00000603
    );
  blk00000001_blk0000044c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000730,
      Q => blk00000001_sig00000604
    );
  blk00000001_blk0000044b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000731,
      Q => blk00000001_sig00000605
    );
  blk00000001_blk0000044a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000732,
      Q => blk00000001_sig00000606
    );
  blk00000001_blk00000449 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000733,
      Q => blk00000001_sig00000607
    );
  blk00000001_blk00000448 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000734,
      Q => blk00000001_sig00000608
    );
  blk00000001_blk00000447 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000735,
      Q => blk00000001_sig00000609
    );
  blk00000001_blk00000446 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000736,
      Q => blk00000001_sig0000060a
    );
  blk00000001_blk00000445 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000737,
      Q => blk00000001_sig0000060b
    );
  blk00000001_blk00000444 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000738,
      Q => blk00000001_sig0000060c
    );
  blk00000001_blk00000443 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000739,
      Q => blk00000001_sig0000060d
    );
  blk00000001_blk00000442 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073a,
      Q => blk00000001_sig0000060e
    );
  blk00000001_blk00000441 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073b,
      Q => blk00000001_sig0000060f
    );
  blk00000001_blk00000440 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073c,
      Q => blk00000001_sig00000610
    );
  blk00000001_blk0000043f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073d,
      Q => blk00000001_sig00000611
    );
  blk00000001_blk0000043e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073e,
      Q => blk00000001_sig00000612
    );
  blk00000001_blk0000043d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000073f,
      Q => blk00000001_sig00000613
    );
  blk00000001_blk0000043c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000740,
      Q => blk00000001_sig00000614
    );
  blk00000001_blk0000043b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000741,
      Q => blk00000001_sig00000615
    );
  blk00000001_blk0000043a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071a,
      Q => blk00000001_sig000005ee
    );
  blk00000001_blk00000439 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071b,
      Q => blk00000001_sig000005ef
    );
  blk00000001_blk00000438 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071c,
      Q => blk00000001_sig000005f0
    );
  blk00000001_blk00000437 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071d,
      Q => blk00000001_sig000005f1
    );
  blk00000001_blk00000436 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071e,
      Q => blk00000001_sig000005f2
    );
  blk00000001_blk00000435 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000071f,
      Q => blk00000001_sig000005f3
    );
  blk00000001_blk00000434 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000720,
      Q => blk00000001_sig000005f4
    );
  blk00000001_blk00000433 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000721,
      Q => blk00000001_sig000005f5
    );
  blk00000001_blk00000432 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000722,
      Q => blk00000001_sig000005f6
    );
  blk00000001_blk00000431 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000723,
      Q => blk00000001_sig000005f7
    );
  blk00000001_blk00000430 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000724,
      Q => blk00000001_sig000005f8
    );
  blk00000001_blk0000042f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000725,
      Q => blk00000001_sig000005f9
    );
  blk00000001_blk0000042e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000726,
      Q => blk00000001_sig000005fa
    );
  blk00000001_blk0000042d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000727,
      Q => blk00000001_sig000005fb
    );
  blk00000001_blk0000042c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000728,
      Q => blk00000001_sig000005fc
    );
  blk00000001_blk0000042b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000729,
      Q => blk00000001_sig000005fd
    );
  blk00000001_blk0000042a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072a,
      Q => blk00000001_sig000005fe
    );
  blk00000001_blk00000429 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072b,
      Q => blk00000001_sig000005ff
    );
  blk00000001_blk00000428 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072c,
      Q => blk00000001_sig00000600
    );
  blk00000001_blk00000427 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000072d,
      Q => blk00000001_sig00000601
    );
  blk00000001_blk00000426 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000706,
      Q => blk00000001_sig000005da
    );
  blk00000001_blk00000425 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000707,
      Q => blk00000001_sig000005db
    );
  blk00000001_blk00000424 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000708,
      Q => blk00000001_sig000005dc
    );
  blk00000001_blk00000423 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000709,
      Q => blk00000001_sig000005dd
    );
  blk00000001_blk00000422 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070a,
      Q => blk00000001_sig000005de
    );
  blk00000001_blk00000421 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070b,
      Q => blk00000001_sig000005df
    );
  blk00000001_blk00000420 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070c,
      Q => blk00000001_sig000005e0
    );
  blk00000001_blk0000041f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070d,
      Q => blk00000001_sig000005e1
    );
  blk00000001_blk0000041e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070e,
      Q => blk00000001_sig000005e2
    );
  blk00000001_blk0000041d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000070f,
      Q => blk00000001_sig000005e3
    );
  blk00000001_blk0000041c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000710,
      Q => blk00000001_sig000005e4
    );
  blk00000001_blk0000041b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000711,
      Q => blk00000001_sig000005e5
    );
  blk00000001_blk0000041a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000712,
      Q => blk00000001_sig000005e6
    );
  blk00000001_blk00000419 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000713,
      Q => blk00000001_sig000005e7
    );
  blk00000001_blk00000418 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000714,
      Q => blk00000001_sig000005e8
    );
  blk00000001_blk00000417 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000715,
      Q => blk00000001_sig000005e9
    );
  blk00000001_blk00000416 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000716,
      Q => blk00000001_sig000005ea
    );
  blk00000001_blk00000415 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000717,
      Q => blk00000001_sig000005eb
    );
  blk00000001_blk00000414 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000718,
      Q => blk00000001_sig000005ec
    );
  blk00000001_blk00000413 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000719,
      Q => blk00000001_sig000005ed
    );
  blk00000001_blk00000412 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f2,
      Q => blk00000001_sig000005c6
    );
  blk00000001_blk00000411 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f3,
      Q => blk00000001_sig000005c7
    );
  blk00000001_blk00000410 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f4,
      Q => blk00000001_sig000005c8
    );
  blk00000001_blk0000040f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f5,
      Q => blk00000001_sig000005c9
    );
  blk00000001_blk0000040e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f6,
      Q => blk00000001_sig000005ca
    );
  blk00000001_blk0000040d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f7,
      Q => blk00000001_sig000005cb
    );
  blk00000001_blk0000040c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f8,
      Q => blk00000001_sig000005cc
    );
  blk00000001_blk0000040b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f9,
      Q => blk00000001_sig000005cd
    );
  blk00000001_blk0000040a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006fa,
      Q => blk00000001_sig000005ce
    );
  blk00000001_blk00000409 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006fb,
      Q => blk00000001_sig000005cf
    );
  blk00000001_blk00000408 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006fc,
      Q => blk00000001_sig000005d0
    );
  blk00000001_blk00000407 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006fd,
      Q => blk00000001_sig000005d1
    );
  blk00000001_blk00000406 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006fe,
      Q => blk00000001_sig000005d2
    );
  blk00000001_blk00000405 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ff,
      Q => blk00000001_sig000005d3
    );
  blk00000001_blk00000404 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000700,
      Q => blk00000001_sig000005d4
    );
  blk00000001_blk00000403 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000701,
      Q => blk00000001_sig000005d5
    );
  blk00000001_blk00000402 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000702,
      Q => blk00000001_sig000005d6
    );
  blk00000001_blk00000401 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000703,
      Q => blk00000001_sig000005d7
    );
  blk00000001_blk00000400 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000704,
      Q => blk00000001_sig000005d8
    );
  blk00000001_blk000003ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000705,
      Q => blk00000001_sig000005d9
    );
  blk00000001_blk000003fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006de,
      Q => blk00000001_sig000005b2
    );
  blk00000001_blk000003fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006df,
      Q => blk00000001_sig000005b3
    );
  blk00000001_blk000003fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e0,
      Q => blk00000001_sig000005b4
    );
  blk00000001_blk000003fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e1,
      Q => blk00000001_sig000005b5
    );
  blk00000001_blk000003fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e2,
      Q => blk00000001_sig000005b6
    );
  blk00000001_blk000003f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e3,
      Q => blk00000001_sig000005b7
    );
  blk00000001_blk000003f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e4,
      Q => blk00000001_sig000005b8
    );
  blk00000001_blk000003f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e5,
      Q => blk00000001_sig000005b9
    );
  blk00000001_blk000003f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e6,
      Q => blk00000001_sig000005ba
    );
  blk00000001_blk000003f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e7,
      Q => blk00000001_sig000005bb
    );
  blk00000001_blk000003f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e8,
      Q => blk00000001_sig000005bc
    );
  blk00000001_blk000003f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006e9,
      Q => blk00000001_sig000005bd
    );
  blk00000001_blk000003f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ea,
      Q => blk00000001_sig000005be
    );
  blk00000001_blk000003f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006eb,
      Q => blk00000001_sig000005bf
    );
  blk00000001_blk000003f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ec,
      Q => blk00000001_sig000005c0
    );
  blk00000001_blk000003ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ed,
      Q => blk00000001_sig000005c1
    );
  blk00000001_blk000003ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ee,
      Q => blk00000001_sig000005c2
    );
  blk00000001_blk000003ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ef,
      Q => blk00000001_sig000005c3
    );
  blk00000001_blk000003ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f0,
      Q => blk00000001_sig000005c4
    );
  blk00000001_blk000003eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006f1,
      Q => blk00000001_sig000005c5
    );
  blk00000001_blk000003ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000742,
      Q => blk00000001_sig000004ee
    );
  blk00000001_blk000003e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000743,
      Q => blk00000001_sig000004ef
    );
  blk00000001_blk000003e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000744,
      Q => blk00000001_sig000004f0
    );
  blk00000001_blk000003e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000745,
      Q => blk00000001_sig000004f1
    );
  blk00000001_blk000003e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000746,
      Q => blk00000001_sig000004f2
    );
  blk00000001_blk000003e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000747,
      Q => blk00000001_sig000004f3
    );
  blk00000001_blk000003e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000748,
      Q => blk00000001_sig000004f4
    );
  blk00000001_blk000003e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000749,
      Q => blk00000001_sig000004f5
    );
  blk00000001_blk000003e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074a,
      Q => blk00000001_sig000004f6
    );
  blk00000001_blk000003e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074b,
      Q => blk00000001_sig000004f7
    );
  blk00000001_blk000003e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074c,
      Q => blk00000001_sig000004f8
    );
  blk00000001_blk000003df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074d,
      Q => blk00000001_sig000004f9
    );
  blk00000001_blk000003de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074e,
      Q => blk00000001_sig000004fa
    );
  blk00000001_blk000003dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000074f,
      Q => blk00000001_sig000004fb
    );
  blk00000001_blk000003dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000750,
      Q => blk00000001_sig000004fc
    );
  blk00000001_blk000003db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000751,
      Q => blk00000001_sig000004fd
    );
  blk00000001_blk000003da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000752,
      Q => blk00000001_sig000004fe
    );
  blk00000001_blk000003d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000753,
      Q => blk00000001_sig000004ff
    );
  blk00000001_blk000003d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000754,
      Q => blk00000001_sig00000500
    );
  blk00000001_blk000003d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000755,
      Q => blk00000001_sig00000501
    );
  blk00000001_blk000003d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069a,
      Q => blk00000001_sig00000586
    );
  blk00000001_blk000003d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069b,
      Q => blk00000001_sig00000587
    );
  blk00000001_blk000003d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069c,
      Q => blk00000001_sig00000588
    );
  blk00000001_blk000003d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069d,
      Q => blk00000001_sig00000589
    );
  blk00000001_blk000003d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069e,
      Q => blk00000001_sig0000058a
    );
  blk00000001_blk000003d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000069f,
      Q => blk00000001_sig0000058b
    );
  blk00000001_blk000003d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a0,
      Q => blk00000001_sig0000058c
    );
  blk00000001_blk000003cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a1,
      Q => blk00000001_sig0000058d
    );
  blk00000001_blk000003ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a2,
      Q => blk00000001_sig0000058e
    );
  blk00000001_blk000003cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a3,
      Q => blk00000001_sig0000058f
    );
  blk00000001_blk000003cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a4,
      Q => blk00000001_sig00000590
    );
  blk00000001_blk000003cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a5,
      Q => blk00000001_sig00000591
    );
  blk00000001_blk000003ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a6,
      Q => blk00000001_sig00000592
    );
  blk00000001_blk000003c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a7,
      Q => blk00000001_sig00000593
    );
  blk00000001_blk000003c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a8,
      Q => blk00000001_sig00000594
    );
  blk00000001_blk000003c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006a9,
      Q => blk00000001_sig00000595
    );
  blk00000001_blk000003c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006aa,
      Q => blk00000001_sig00000596
    );
  blk00000001_blk000003c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ab,
      Q => blk00000001_sig00000597
    );
  blk00000001_blk000003c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ac,
      Q => blk00000001_sig00000598
    );
  blk00000001_blk000003c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ad,
      Q => blk00000001_sig00000599
    );
  blk00000001_blk000003c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ae,
      Q => blk00000001_sig0000059a
    );
  blk00000001_blk000003c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006af,
      Q => blk00000001_sig0000059b
    );
  blk00000001_blk000003c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b0,
      Q => blk00000001_sig0000059c
    );
  blk00000001_blk000003bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b1,
      Q => blk00000001_sig0000059d
    );
  blk00000001_blk000003be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b2,
      Q => blk00000001_sig0000059e
    );
  blk00000001_blk000003bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b3,
      Q => blk00000001_sig0000059f
    );
  blk00000001_blk000003bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b4,
      Q => blk00000001_sig000005a0
    );
  blk00000001_blk000003bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b5,
      Q => blk00000001_sig000005a1
    );
  blk00000001_blk000003ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b6,
      Q => blk00000001_sig000005a2
    );
  blk00000001_blk000003b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b7,
      Q => blk00000001_sig000005a3
    );
  blk00000001_blk000003b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b8,
      Q => blk00000001_sig000005a4
    );
  blk00000001_blk000003b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006b9,
      Q => blk00000001_sig000005a5
    );
  blk00000001_blk000003b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006ba,
      Q => blk00000001_sig000005a6
    );
  blk00000001_blk000003b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006bb,
      Q => blk00000001_sig000005a7
    );
  blk00000001_blk000003b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006bc,
      Q => blk00000001_sig000005a8
    );
  blk00000001_blk000003b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006bd,
      Q => blk00000001_sig000005a9
    );
  blk00000001_blk000003b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006be,
      Q => blk00000001_sig000005aa
    );
  blk00000001_blk000003b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006bf,
      Q => blk00000001_sig000005ab
    );
  blk00000001_blk000003b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c0,
      Q => blk00000001_sig000005ac
    );
  blk00000001_blk000003af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c1,
      Q => blk00000001_sig000005ad
    );
  blk00000001_blk000003ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c2,
      Q => blk00000001_sig000005ae
    );
  blk00000001_blk000003ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c3,
      Q => blk00000001_sig000005af
    );
  blk00000001_blk000003ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c4,
      Q => blk00000001_sig000005b0
    );
  blk00000001_blk000003ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000006c5,
      Q => blk00000001_sig000005b1
    );
  blk00000001_blk000003aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000658,
      Q => blk00000001_sig00000570
    );
  blk00000001_blk000003a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000659,
      Q => blk00000001_sig00000571
    );
  blk00000001_blk000003a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065a,
      Q => blk00000001_sig00000572
    );
  blk00000001_blk000003a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065b,
      Q => blk00000001_sig00000573
    );
  blk00000001_blk000003a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065c,
      Q => blk00000001_sig00000574
    );
  blk00000001_blk000003a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065d,
      Q => blk00000001_sig00000575
    );
  blk00000001_blk000003a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065e,
      Q => blk00000001_sig00000576
    );
  blk00000001_blk000003a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000065f,
      Q => blk00000001_sig00000577
    );
  blk00000001_blk000003a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000660,
      Q => blk00000001_sig00000578
    );
  blk00000001_blk000003a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000661,
      Q => blk00000001_sig00000579
    );
  blk00000001_blk000003a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000662,
      Q => blk00000001_sig0000057a
    );
  blk00000001_blk0000039f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000663,
      Q => blk00000001_sig0000057b
    );
  blk00000001_blk0000039e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000664,
      Q => blk00000001_sig0000057c
    );
  blk00000001_blk0000039d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000665,
      Q => blk00000001_sig0000057d
    );
  blk00000001_blk0000039c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000666,
      Q => blk00000001_sig0000057e
    );
  blk00000001_blk0000039b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000667,
      Q => blk00000001_sig0000057f
    );
  blk00000001_blk0000039a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000668,
      Q => blk00000001_sig00000580
    );
  blk00000001_blk00000399 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000669,
      Q => blk00000001_sig00000581
    );
  blk00000001_blk00000398 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066a,
      Q => blk00000001_sig00000582
    );
  blk00000001_blk00000397 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066b,
      Q => blk00000001_sig00000583
    );
  blk00000001_blk00000396 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066c,
      Q => blk00000001_sig00000584
    );
  blk00000001_blk00000395 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066d,
      Q => blk00000001_sig00000585
    );
  blk00000001_blk00000394 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000642,
      Q => blk00000001_sig0000055a
    );
  blk00000001_blk00000393 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000643,
      Q => blk00000001_sig0000055b
    );
  blk00000001_blk00000392 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000644,
      Q => blk00000001_sig0000055c
    );
  blk00000001_blk00000391 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000645,
      Q => blk00000001_sig0000055d
    );
  blk00000001_blk00000390 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000646,
      Q => blk00000001_sig0000055e
    );
  blk00000001_blk0000038f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000647,
      Q => blk00000001_sig0000055f
    );
  blk00000001_blk0000038e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000648,
      Q => blk00000001_sig00000560
    );
  blk00000001_blk0000038d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000649,
      Q => blk00000001_sig00000561
    );
  blk00000001_blk0000038c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064a,
      Q => blk00000001_sig00000562
    );
  blk00000001_blk0000038b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064b,
      Q => blk00000001_sig00000563
    );
  blk00000001_blk0000038a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064c,
      Q => blk00000001_sig00000564
    );
  blk00000001_blk00000389 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064d,
      Q => blk00000001_sig00000565
    );
  blk00000001_blk00000388 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064e,
      Q => blk00000001_sig00000566
    );
  blk00000001_blk00000387 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000064f,
      Q => blk00000001_sig00000567
    );
  blk00000001_blk00000386 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000650,
      Q => blk00000001_sig00000568
    );
  blk00000001_blk00000385 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000651,
      Q => blk00000001_sig00000569
    );
  blk00000001_blk00000384 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000652,
      Q => blk00000001_sig0000056a
    );
  blk00000001_blk00000383 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000653,
      Q => blk00000001_sig0000056b
    );
  blk00000001_blk00000382 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000654,
      Q => blk00000001_sig0000056c
    );
  blk00000001_blk00000381 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000655,
      Q => blk00000001_sig0000056d
    );
  blk00000001_blk00000380 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000656,
      Q => blk00000001_sig0000056e
    );
  blk00000001_blk0000037f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000657,
      Q => blk00000001_sig0000056f
    );
  blk00000001_blk0000037e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000684,
      Q => blk00000001_sig00000544
    );
  blk00000001_blk0000037d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000685,
      Q => blk00000001_sig00000545
    );
  blk00000001_blk0000037c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000686,
      Q => blk00000001_sig00000546
    );
  blk00000001_blk0000037b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000687,
      Q => blk00000001_sig00000547
    );
  blk00000001_blk0000037a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000688,
      Q => blk00000001_sig00000548
    );
  blk00000001_blk00000379 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000689,
      Q => blk00000001_sig00000549
    );
  blk00000001_blk00000378 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068a,
      Q => blk00000001_sig0000054a
    );
  blk00000001_blk00000377 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068b,
      Q => blk00000001_sig0000054b
    );
  blk00000001_blk00000376 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068c,
      Q => blk00000001_sig0000054c
    );
  blk00000001_blk00000375 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068d,
      Q => blk00000001_sig0000054d
    );
  blk00000001_blk00000374 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068e,
      Q => blk00000001_sig0000054e
    );
  blk00000001_blk00000373 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000068f,
      Q => blk00000001_sig0000054f
    );
  blk00000001_blk00000372 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000690,
      Q => blk00000001_sig00000550
    );
  blk00000001_blk00000371 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000691,
      Q => blk00000001_sig00000551
    );
  blk00000001_blk00000370 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000692,
      Q => blk00000001_sig00000552
    );
  blk00000001_blk0000036f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000693,
      Q => blk00000001_sig00000553
    );
  blk00000001_blk0000036e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000694,
      Q => blk00000001_sig00000554
    );
  blk00000001_blk0000036d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000695,
      Q => blk00000001_sig00000555
    );
  blk00000001_blk0000036c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000696,
      Q => blk00000001_sig00000556
    );
  blk00000001_blk0000036b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000697,
      Q => blk00000001_sig00000557
    );
  blk00000001_blk0000036a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000698,
      Q => blk00000001_sig00000558
    );
  blk00000001_blk00000369 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000699,
      Q => blk00000001_sig00000559
    );
  blk00000001_blk00000368 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066e,
      Q => blk00000001_sig0000052e
    );
  blk00000001_blk00000367 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000066f,
      Q => blk00000001_sig0000052f
    );
  blk00000001_blk00000366 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000670,
      Q => blk00000001_sig00000530
    );
  blk00000001_blk00000365 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000671,
      Q => blk00000001_sig00000531
    );
  blk00000001_blk00000364 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000672,
      Q => blk00000001_sig00000532
    );
  blk00000001_blk00000363 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000673,
      Q => blk00000001_sig00000533
    );
  blk00000001_blk00000362 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000674,
      Q => blk00000001_sig00000534
    );
  blk00000001_blk00000361 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000675,
      Q => blk00000001_sig00000535
    );
  blk00000001_blk00000360 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000676,
      Q => blk00000001_sig00000536
    );
  blk00000001_blk0000035f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000677,
      Q => blk00000001_sig00000537
    );
  blk00000001_blk0000035e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000678,
      Q => blk00000001_sig00000538
    );
  blk00000001_blk0000035d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000679,
      Q => blk00000001_sig00000539
    );
  blk00000001_blk0000035c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067a,
      Q => blk00000001_sig0000053a
    );
  blk00000001_blk0000035b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067b,
      Q => blk00000001_sig0000053b
    );
  blk00000001_blk0000035a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067c,
      Q => blk00000001_sig0000053c
    );
  blk00000001_blk00000359 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067d,
      Q => blk00000001_sig0000053d
    );
  blk00000001_blk00000358 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067e,
      Q => blk00000001_sig0000053e
    );
  blk00000001_blk00000357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000067f,
      Q => blk00000001_sig0000053f
    );
  blk00000001_blk00000356 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000680,
      Q => blk00000001_sig00000540
    );
  blk00000001_blk00000355 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000681,
      Q => blk00000001_sig00000541
    );
  blk00000001_blk00000354 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000682,
      Q => blk00000001_sig00000542
    );
  blk00000001_blk00000353 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000683,
      Q => blk00000001_sig00000543
    );
  blk00000001_blk00000352 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062c,
      Q => blk00000001_sig00000518
    );
  blk00000001_blk00000351 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062d,
      Q => blk00000001_sig00000519
    );
  blk00000001_blk00000350 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062e,
      Q => blk00000001_sig0000051a
    );
  blk00000001_blk0000034f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062f,
      Q => blk00000001_sig0000051b
    );
  blk00000001_blk0000034e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000630,
      Q => blk00000001_sig0000051c
    );
  blk00000001_blk0000034d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000631,
      Q => blk00000001_sig0000051d
    );
  blk00000001_blk0000034c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000632,
      Q => blk00000001_sig0000051e
    );
  blk00000001_blk0000034b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000633,
      Q => blk00000001_sig0000051f
    );
  blk00000001_blk0000034a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000634,
      Q => blk00000001_sig00000520
    );
  blk00000001_blk00000349 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000635,
      Q => blk00000001_sig00000521
    );
  blk00000001_blk00000348 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000636,
      Q => blk00000001_sig00000522
    );
  blk00000001_blk00000347 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000637,
      Q => blk00000001_sig00000523
    );
  blk00000001_blk00000346 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000638,
      Q => blk00000001_sig00000524
    );
  blk00000001_blk00000345 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000639,
      Q => blk00000001_sig00000525
    );
  blk00000001_blk00000344 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063a,
      Q => blk00000001_sig00000526
    );
  blk00000001_blk00000343 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063b,
      Q => blk00000001_sig00000527
    );
  blk00000001_blk00000342 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063c,
      Q => blk00000001_sig00000528
    );
  blk00000001_blk00000341 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063d,
      Q => blk00000001_sig00000529
    );
  blk00000001_blk00000340 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063e,
      Q => blk00000001_sig0000052a
    );
  blk00000001_blk0000033f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000063f,
      Q => blk00000001_sig0000052b
    );
  blk00000001_blk0000033e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000640,
      Q => blk00000001_sig0000052c
    );
  blk00000001_blk0000033d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000641,
      Q => blk00000001_sig0000052d
    );
  blk00000001_blk0000033c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000616,
      Q => blk00000001_sig00000502
    );
  blk00000001_blk0000033b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000617,
      Q => blk00000001_sig00000503
    );
  blk00000001_blk0000033a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000618,
      Q => blk00000001_sig00000504
    );
  blk00000001_blk00000339 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000619,
      Q => blk00000001_sig00000505
    );
  blk00000001_blk00000338 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061a,
      Q => blk00000001_sig00000506
    );
  blk00000001_blk00000337 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061b,
      Q => blk00000001_sig00000507
    );
  blk00000001_blk00000336 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061c,
      Q => blk00000001_sig00000508
    );
  blk00000001_blk00000335 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061d,
      Q => blk00000001_sig00000509
    );
  blk00000001_blk00000334 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061e,
      Q => blk00000001_sig0000050a
    );
  blk00000001_blk00000333 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000061f,
      Q => blk00000001_sig0000050b
    );
  blk00000001_blk00000332 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000620,
      Q => blk00000001_sig0000050c
    );
  blk00000001_blk00000331 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000621,
      Q => blk00000001_sig0000050d
    );
  blk00000001_blk00000330 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000622,
      Q => blk00000001_sig0000050e
    );
  blk00000001_blk0000032f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000623,
      Q => blk00000001_sig0000050f
    );
  blk00000001_blk0000032e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000624,
      Q => blk00000001_sig00000510
    );
  blk00000001_blk0000032d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000625,
      Q => blk00000001_sig00000511
    );
  blk00000001_blk0000032c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000626,
      Q => blk00000001_sig00000512
    );
  blk00000001_blk0000032b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000627,
      Q => blk00000001_sig00000513
    );
  blk00000001_blk0000032a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000628,
      Q => blk00000001_sig00000514
    );
  blk00000001_blk00000329 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000629,
      Q => blk00000001_sig00000515
    );
  blk00000001_blk00000328 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062a,
      Q => blk00000001_sig00000516
    );
  blk00000001_blk00000327 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000062b,
      Q => blk00000001_sig00000517
    );
  blk00000001_blk00000326 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004ed,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000009b
    );
  blk00000001_blk00000325 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004ec,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000009c
    );
  blk00000001_blk00000324 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004eb,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000009d
    );
  blk00000001_blk00000323 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004ea,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000009e
    );
  blk00000001_blk00000322 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000009f
    );
  blk00000001_blk00000321 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a0
    );
  blk00000001_blk00000320 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a1
    );
  blk00000001_blk0000031f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a2
    );
  blk00000001_blk0000031e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a3
    );
  blk00000001_blk0000031d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a4
    );
  blk00000001_blk0000031c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a5
    );
  blk00000001_blk0000031b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a6
    );
  blk00000001_blk0000031a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a7
    );
  blk00000001_blk00000319 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004e0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a8
    );
  blk00000001_blk00000318 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004df,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000a9
    );
  blk00000001_blk00000317 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004de,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000aa
    );
  blk00000001_blk00000316 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000200,
      I1 => blk00000001_sig00000220,
      I2 => blk00000001_sig00000240,
      I3 => blk00000001_sig00000260,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004ed
    );
  blk00000001_blk00000315 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ff,
      I1 => blk00000001_sig0000021f,
      I2 => blk00000001_sig0000023f,
      I3 => blk00000001_sig0000025f,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004ec
    );
  blk00000001_blk00000314 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fe,
      I1 => blk00000001_sig0000021e,
      I2 => blk00000001_sig0000023e,
      I3 => blk00000001_sig0000025e,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004eb
    );
  blk00000001_blk00000313 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fd,
      I1 => blk00000001_sig0000021d,
      I2 => blk00000001_sig0000023d,
      I3 => blk00000001_sig0000025d,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004ea
    );
  blk00000001_blk00000312 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fc,
      I1 => blk00000001_sig0000021c,
      I2 => blk00000001_sig0000023c,
      I3 => blk00000001_sig0000025c,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e9
    );
  blk00000001_blk00000311 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fb,
      I1 => blk00000001_sig0000021b,
      I2 => blk00000001_sig0000023b,
      I3 => blk00000001_sig0000025b,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e8
    );
  blk00000001_blk00000310 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fa,
      I1 => blk00000001_sig0000021a,
      I2 => blk00000001_sig0000023a,
      I3 => blk00000001_sig0000025a,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e7
    );
  blk00000001_blk0000030f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f9,
      I1 => blk00000001_sig00000219,
      I2 => blk00000001_sig00000239,
      I3 => blk00000001_sig00000259,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e6
    );
  blk00000001_blk0000030e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f8,
      I1 => blk00000001_sig00000218,
      I2 => blk00000001_sig00000238,
      I3 => blk00000001_sig00000258,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e5
    );
  blk00000001_blk0000030d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f7,
      I1 => blk00000001_sig00000217,
      I2 => blk00000001_sig00000237,
      I3 => blk00000001_sig00000257,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e4
    );
  blk00000001_blk0000030c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f6,
      I1 => blk00000001_sig00000216,
      I2 => blk00000001_sig00000236,
      I3 => blk00000001_sig00000256,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e3
    );
  blk00000001_blk0000030b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f5,
      I1 => blk00000001_sig00000215,
      I2 => blk00000001_sig00000235,
      I3 => blk00000001_sig00000255,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e2
    );
  blk00000001_blk0000030a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f4,
      I1 => blk00000001_sig00000214,
      I2 => blk00000001_sig00000234,
      I3 => blk00000001_sig00000254,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e1
    );
  blk00000001_blk00000309 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f3,
      I1 => blk00000001_sig00000213,
      I2 => blk00000001_sig00000233,
      I3 => blk00000001_sig00000253,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004e0
    );
  blk00000001_blk00000308 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f2,
      I1 => blk00000001_sig00000212,
      I2 => blk00000001_sig00000232,
      I3 => blk00000001_sig00000252,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004df
    );
  blk00000001_blk00000307 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f1,
      I1 => blk00000001_sig00000211,
      I2 => blk00000001_sig00000231,
      I3 => blk00000001_sig00000251,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004de
    );
  blk00000001_blk00000306 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004dd,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000ab
    );
  blk00000001_blk00000305 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004dc,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000ac
    );
  blk00000001_blk00000304 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004db,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000ad
    );
  blk00000001_blk00000303 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004da,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000ae
    );
  blk00000001_blk00000302 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d9,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000af
    );
  blk00000001_blk00000301 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d8,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b0
    );
  blk00000001_blk00000300 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d7,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b1
    );
  blk00000001_blk000002ff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d6,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b2
    );
  blk00000001_blk000002fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d5,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b3
    );
  blk00000001_blk000002fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d4,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b4
    );
  blk00000001_blk000002fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d3,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b5
    );
  blk00000001_blk000002fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d2,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b6
    );
  blk00000001_blk000002fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d1,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b7
    );
  blk00000001_blk000002f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004d0,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b8
    );
  blk00000001_blk000002f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004cf,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000b9
    );
  blk00000001_blk000002f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000004ce,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig000000ba
    );
  blk00000001_blk000002f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f0,
      I1 => blk00000001_sig00000210,
      I2 => blk00000001_sig00000230,
      I3 => blk00000001_sig00000250,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004dd
    );
  blk00000001_blk000002f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ef,
      I1 => blk00000001_sig0000020f,
      I2 => blk00000001_sig0000022f,
      I3 => blk00000001_sig0000024f,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004dc
    );
  blk00000001_blk000002f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ee,
      I1 => blk00000001_sig0000020e,
      I2 => blk00000001_sig0000022e,
      I3 => blk00000001_sig0000024e,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004db
    );
  blk00000001_blk000002f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ed,
      I1 => blk00000001_sig0000020d,
      I2 => blk00000001_sig0000022d,
      I3 => blk00000001_sig0000024d,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004da
    );
  blk00000001_blk000002f2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ec,
      I1 => blk00000001_sig0000020c,
      I2 => blk00000001_sig0000022c,
      I3 => blk00000001_sig0000024c,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d9
    );
  blk00000001_blk000002f1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001eb,
      I1 => blk00000001_sig0000020b,
      I2 => blk00000001_sig0000022b,
      I3 => blk00000001_sig0000024b,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d8
    );
  blk00000001_blk000002f0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ea,
      I1 => blk00000001_sig0000020a,
      I2 => blk00000001_sig0000022a,
      I3 => blk00000001_sig0000024a,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d7
    );
  blk00000001_blk000002ef : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e9,
      I1 => blk00000001_sig00000209,
      I2 => blk00000001_sig00000229,
      I3 => blk00000001_sig00000249,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d6
    );
  blk00000001_blk000002ee : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e8,
      I1 => blk00000001_sig00000208,
      I2 => blk00000001_sig00000228,
      I3 => blk00000001_sig00000248,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d5
    );
  blk00000001_blk000002ed : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e7,
      I1 => blk00000001_sig00000207,
      I2 => blk00000001_sig00000227,
      I3 => blk00000001_sig00000247,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d4
    );
  blk00000001_blk000002ec : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e6,
      I1 => blk00000001_sig00000206,
      I2 => blk00000001_sig00000226,
      I3 => blk00000001_sig00000246,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d3
    );
  blk00000001_blk000002eb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e5,
      I1 => blk00000001_sig00000205,
      I2 => blk00000001_sig00000225,
      I3 => blk00000001_sig00000245,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d2
    );
  blk00000001_blk000002ea : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e4,
      I1 => blk00000001_sig00000204,
      I2 => blk00000001_sig00000224,
      I3 => blk00000001_sig00000244,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d1
    );
  blk00000001_blk000002e9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e3,
      I1 => blk00000001_sig00000203,
      I2 => blk00000001_sig00000223,
      I3 => blk00000001_sig00000243,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004d0
    );
  blk00000001_blk000002e8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e2,
      I1 => blk00000001_sig00000202,
      I2 => blk00000001_sig00000222,
      I3 => blk00000001_sig00000242,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004cf
    );
  blk00000001_blk000002e7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e1,
      I1 => blk00000001_sig00000201,
      I2 => blk00000001_sig00000221,
      I3 => blk00000001_sig00000241,
      I4 => blk00000001_sig000001b3,
      I5 => blk00000001_sig000001b4,
      O => blk00000001_sig000004ce
    );
  blk00000001_blk000002e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004cd,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f7
    );
  blk00000001_blk000002e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004cc,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f6
    );
  blk00000001_blk000002e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004cb,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f5
    );
  blk00000001_blk000002e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ca,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f4
    );
  blk00000001_blk000002e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c9,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f3
    );
  blk00000001_blk000002e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c8,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f2
    );
  blk00000001_blk000002e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c7,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f1
    );
  blk00000001_blk000002df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c6,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f0
    );
  blk00000001_blk000002de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c5,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ef
    );
  blk00000001_blk000002dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c4,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ee
    );
  blk00000001_blk000002dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c3,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ed
    );
  blk00000001_blk000002db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c2,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ec
    );
  blk00000001_blk000002da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c1,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003eb
    );
  blk00000001_blk000002d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004c0,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ea
    );
  blk00000001_blk000002d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004bf,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003e9
    );
  blk00000001_blk000002d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004be,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003e8
    );
  blk00000001_blk000002d6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f0,
      I1 => blk00000001_sig00000210,
      I2 => blk00000001_sig00000230,
      I3 => blk00000001_sig00000250,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004cd
    );
  blk00000001_blk000002d5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ef,
      I1 => blk00000001_sig0000020f,
      I2 => blk00000001_sig0000022f,
      I3 => blk00000001_sig0000024f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004cc
    );
  blk00000001_blk000002d4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ee,
      I1 => blk00000001_sig0000020e,
      I2 => blk00000001_sig0000022e,
      I3 => blk00000001_sig0000024e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004cb
    );
  blk00000001_blk000002d3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ed,
      I1 => blk00000001_sig0000020d,
      I2 => blk00000001_sig0000022d,
      I3 => blk00000001_sig0000024d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ca
    );
  blk00000001_blk000002d2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ec,
      I1 => blk00000001_sig0000020c,
      I2 => blk00000001_sig0000022c,
      I3 => blk00000001_sig0000024c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c9
    );
  blk00000001_blk000002d1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001eb,
      I1 => blk00000001_sig0000020b,
      I2 => blk00000001_sig0000022b,
      I3 => blk00000001_sig0000024b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c8
    );
  blk00000001_blk000002d0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ea,
      I1 => blk00000001_sig0000020a,
      I2 => blk00000001_sig0000022a,
      I3 => blk00000001_sig0000024a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c7
    );
  blk00000001_blk000002cf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e9,
      I1 => blk00000001_sig00000209,
      I2 => blk00000001_sig00000229,
      I3 => blk00000001_sig00000249,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c6
    );
  blk00000001_blk000002ce : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e8,
      I1 => blk00000001_sig00000208,
      I2 => blk00000001_sig00000228,
      I3 => blk00000001_sig00000248,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c5
    );
  blk00000001_blk000002cd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e7,
      I1 => blk00000001_sig00000207,
      I2 => blk00000001_sig00000227,
      I3 => blk00000001_sig00000247,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c4
    );
  blk00000001_blk000002cc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e6,
      I1 => blk00000001_sig00000206,
      I2 => blk00000001_sig00000226,
      I3 => blk00000001_sig00000246,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c3
    );
  blk00000001_blk000002cb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e5,
      I1 => blk00000001_sig00000205,
      I2 => blk00000001_sig00000225,
      I3 => blk00000001_sig00000245,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c2
    );
  blk00000001_blk000002ca : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e4,
      I1 => blk00000001_sig00000204,
      I2 => blk00000001_sig00000224,
      I3 => blk00000001_sig00000244,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c1
    );
  blk00000001_blk000002c9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e3,
      I1 => blk00000001_sig00000203,
      I2 => blk00000001_sig00000223,
      I3 => blk00000001_sig00000243,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004c0
    );
  blk00000001_blk000002c8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e2,
      I1 => blk00000001_sig00000202,
      I2 => blk00000001_sig00000222,
      I3 => blk00000001_sig00000242,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004bf
    );
  blk00000001_blk000002c7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001e1,
      I1 => blk00000001_sig00000201,
      I2 => blk00000001_sig00000221,
      I3 => blk00000001_sig00000241,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004be
    );
  blk00000001_blk000002c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004bd,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d7
    );
  blk00000001_blk000002c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004bc,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d6
    );
  blk00000001_blk000002c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004bb,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d5
    );
  blk00000001_blk000002c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ba,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d4
    );
  blk00000001_blk000002c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b9,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d3
    );
  blk00000001_blk000002c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b8,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d2
    );
  blk00000001_blk000002c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b7,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d1
    );
  blk00000001_blk000002bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b6,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d0
    );
  blk00000001_blk000002be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b5,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007cf
    );
  blk00000001_blk000002bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b4,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007ce
    );
  blk00000001_blk000002bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b3,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007cd
    );
  blk00000001_blk000002bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b2,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007cc
    );
  blk00000001_blk000002ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b1,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007cb
    );
  blk00000001_blk000002b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004b0,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007ca
    );
  blk00000001_blk000002b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004af,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007c9
    );
  blk00000001_blk000002b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ae,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007c8
    );
  blk00000001_blk000002b6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000210,
      I1 => blk00000001_sig00000230,
      I2 => blk00000001_sig00000250,
      I3 => blk00000001_sig000001f0,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004bd
    );
  blk00000001_blk000002b5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020f,
      I1 => blk00000001_sig0000022f,
      I2 => blk00000001_sig0000024f,
      I3 => blk00000001_sig000001ef,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004bc
    );
  blk00000001_blk000002b4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020e,
      I1 => blk00000001_sig0000022e,
      I2 => blk00000001_sig0000024e,
      I3 => blk00000001_sig000001ee,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004bb
    );
  blk00000001_blk000002b3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020d,
      I1 => blk00000001_sig0000022d,
      I2 => blk00000001_sig0000024d,
      I3 => blk00000001_sig000001ed,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ba
    );
  blk00000001_blk000002b2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020c,
      I1 => blk00000001_sig0000022c,
      I2 => blk00000001_sig0000024c,
      I3 => blk00000001_sig000001ec,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b9
    );
  blk00000001_blk000002b1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020b,
      I1 => blk00000001_sig0000022b,
      I2 => blk00000001_sig0000024b,
      I3 => blk00000001_sig000001eb,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b8
    );
  blk00000001_blk000002b0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000020a,
      I1 => blk00000001_sig0000022a,
      I2 => blk00000001_sig0000024a,
      I3 => blk00000001_sig000001ea,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b7
    );
  blk00000001_blk000002af : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000209,
      I1 => blk00000001_sig00000229,
      I2 => blk00000001_sig00000249,
      I3 => blk00000001_sig000001e9,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b6
    );
  blk00000001_blk000002ae : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000208,
      I1 => blk00000001_sig00000228,
      I2 => blk00000001_sig00000248,
      I3 => blk00000001_sig000001e8,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b5
    );
  blk00000001_blk000002ad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000207,
      I1 => blk00000001_sig00000227,
      I2 => blk00000001_sig00000247,
      I3 => blk00000001_sig000001e7,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b4
    );
  blk00000001_blk000002ac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000206,
      I1 => blk00000001_sig00000226,
      I2 => blk00000001_sig00000246,
      I3 => blk00000001_sig000001e6,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b3
    );
  blk00000001_blk000002ab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000205,
      I1 => blk00000001_sig00000225,
      I2 => blk00000001_sig00000245,
      I3 => blk00000001_sig000001e5,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b2
    );
  blk00000001_blk000002aa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000204,
      I1 => blk00000001_sig00000224,
      I2 => blk00000001_sig00000244,
      I3 => blk00000001_sig000001e4,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b1
    );
  blk00000001_blk000002a9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000203,
      I1 => blk00000001_sig00000223,
      I2 => blk00000001_sig00000243,
      I3 => blk00000001_sig000001e3,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004b0
    );
  blk00000001_blk000002a8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000202,
      I1 => blk00000001_sig00000222,
      I2 => blk00000001_sig00000242,
      I3 => blk00000001_sig000001e2,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004af
    );
  blk00000001_blk000002a7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000201,
      I1 => blk00000001_sig00000221,
      I2 => blk00000001_sig00000241,
      I3 => blk00000001_sig000001e1,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ae
    );
  blk00000001_blk000002a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ad,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084a
    );
  blk00000001_blk000002a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ac,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000849
    );
  blk00000001_blk000002a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004ab,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000848
    );
  blk00000001_blk000002a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004aa,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000847
    );
  blk00000001_blk000002a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a9,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000846
    );
  blk00000001_blk000002a1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a8,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000845
    );
  blk00000001_blk000002a0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a7,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000844
    );
  blk00000001_blk0000029f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a6,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000843
    );
  blk00000001_blk0000029e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a5,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000842
    );
  blk00000001_blk0000029d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a4,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000841
    );
  blk00000001_blk0000029c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a3,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000840
    );
  blk00000001_blk0000029b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a2,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000083f
    );
  blk00000001_blk0000029a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a1,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000083e
    );
  blk00000001_blk00000299 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig000004a0,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000083d
    );
  blk00000001_blk00000298 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000083c
    );
  blk00000001_blk00000297 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000083b
    );
  blk00000001_blk00000296 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000230,
      I1 => blk00000001_sig00000250,
      I2 => blk00000001_sig000001f0,
      I3 => blk00000001_sig00000210,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ad
    );
  blk00000001_blk00000295 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022f,
      I1 => blk00000001_sig0000024f,
      I2 => blk00000001_sig000001ef,
      I3 => blk00000001_sig0000020f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ac
    );
  blk00000001_blk00000294 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022e,
      I1 => blk00000001_sig0000024e,
      I2 => blk00000001_sig000001ee,
      I3 => blk00000001_sig0000020e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004ab
    );
  blk00000001_blk00000293 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022d,
      I1 => blk00000001_sig0000024d,
      I2 => blk00000001_sig000001ed,
      I3 => blk00000001_sig0000020d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004aa
    );
  blk00000001_blk00000292 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022c,
      I1 => blk00000001_sig0000024c,
      I2 => blk00000001_sig000001ec,
      I3 => blk00000001_sig0000020c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a9
    );
  blk00000001_blk00000291 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022b,
      I1 => blk00000001_sig0000024b,
      I2 => blk00000001_sig000001eb,
      I3 => blk00000001_sig0000020b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a8
    );
  blk00000001_blk00000290 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000022a,
      I1 => blk00000001_sig0000024a,
      I2 => blk00000001_sig000001ea,
      I3 => blk00000001_sig0000020a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a7
    );
  blk00000001_blk0000028f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000229,
      I1 => blk00000001_sig00000249,
      I2 => blk00000001_sig000001e9,
      I3 => blk00000001_sig00000209,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a6
    );
  blk00000001_blk0000028e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000228,
      I1 => blk00000001_sig00000248,
      I2 => blk00000001_sig000001e8,
      I3 => blk00000001_sig00000208,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a5
    );
  blk00000001_blk0000028d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000227,
      I1 => blk00000001_sig00000247,
      I2 => blk00000001_sig000001e7,
      I3 => blk00000001_sig00000207,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a4
    );
  blk00000001_blk0000028c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000226,
      I1 => blk00000001_sig00000246,
      I2 => blk00000001_sig000001e6,
      I3 => blk00000001_sig00000206,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a3
    );
  blk00000001_blk0000028b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000225,
      I1 => blk00000001_sig00000245,
      I2 => blk00000001_sig000001e5,
      I3 => blk00000001_sig00000205,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a2
    );
  blk00000001_blk0000028a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000224,
      I1 => blk00000001_sig00000244,
      I2 => blk00000001_sig000001e4,
      I3 => blk00000001_sig00000204,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a1
    );
  blk00000001_blk00000289 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000223,
      I1 => blk00000001_sig00000243,
      I2 => blk00000001_sig000001e3,
      I3 => blk00000001_sig00000203,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig000004a0
    );
  blk00000001_blk00000288 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000222,
      I1 => blk00000001_sig00000242,
      I2 => blk00000001_sig000001e2,
      I3 => blk00000001_sig00000202,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049f
    );
  blk00000001_blk00000287 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000221,
      I1 => blk00000001_sig00000241,
      I2 => blk00000001_sig000001e1,
      I3 => blk00000001_sig00000201,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049e
    );
  blk00000001_blk00000286 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049d,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008bf
    );
  blk00000001_blk00000285 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049c,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008be
    );
  blk00000001_blk00000284 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049b,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008bd
    );
  blk00000001_blk00000283 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000049a,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008bc
    );
  blk00000001_blk00000282 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000499,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008bb
    );
  blk00000001_blk00000281 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000498,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008ba
    );
  blk00000001_blk00000280 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000497,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b9
    );
  blk00000001_blk0000027f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000496,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b8
    );
  blk00000001_blk0000027e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000495,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b7
    );
  blk00000001_blk0000027d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000494,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b6
    );
  blk00000001_blk0000027c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000493,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b5
    );
  blk00000001_blk0000027b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000492,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b4
    );
  blk00000001_blk0000027a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000491,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b3
    );
  blk00000001_blk00000279 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000490,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b2
    );
  blk00000001_blk00000278 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b1
    );
  blk00000001_blk00000277 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008b0
    );
  blk00000001_blk00000276 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000250,
      I1 => blk00000001_sig000001f0,
      I2 => blk00000001_sig00000210,
      I3 => blk00000001_sig00000230,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049d
    );
  blk00000001_blk00000275 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024f,
      I1 => blk00000001_sig000001ef,
      I2 => blk00000001_sig0000020f,
      I3 => blk00000001_sig0000022f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049c
    );
  blk00000001_blk00000274 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024e,
      I1 => blk00000001_sig000001ee,
      I2 => blk00000001_sig0000020e,
      I3 => blk00000001_sig0000022e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049b
    );
  blk00000001_blk00000273 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024d,
      I1 => blk00000001_sig000001ed,
      I2 => blk00000001_sig0000020d,
      I3 => blk00000001_sig0000022d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000049a
    );
  blk00000001_blk00000272 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024c,
      I1 => blk00000001_sig000001ec,
      I2 => blk00000001_sig0000020c,
      I3 => blk00000001_sig0000022c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000499
    );
  blk00000001_blk00000271 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024b,
      I1 => blk00000001_sig000001eb,
      I2 => blk00000001_sig0000020b,
      I3 => blk00000001_sig0000022b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000498
    );
  blk00000001_blk00000270 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000024a,
      I1 => blk00000001_sig000001ea,
      I2 => blk00000001_sig0000020a,
      I3 => blk00000001_sig0000022a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000497
    );
  blk00000001_blk0000026f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000249,
      I1 => blk00000001_sig000001e9,
      I2 => blk00000001_sig00000209,
      I3 => blk00000001_sig00000229,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000496
    );
  blk00000001_blk0000026e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000248,
      I1 => blk00000001_sig000001e8,
      I2 => blk00000001_sig00000208,
      I3 => blk00000001_sig00000228,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000495
    );
  blk00000001_blk0000026d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000247,
      I1 => blk00000001_sig000001e7,
      I2 => blk00000001_sig00000207,
      I3 => blk00000001_sig00000227,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000494
    );
  blk00000001_blk0000026c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000246,
      I1 => blk00000001_sig000001e6,
      I2 => blk00000001_sig00000206,
      I3 => blk00000001_sig00000226,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000493
    );
  blk00000001_blk0000026b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000245,
      I1 => blk00000001_sig000001e5,
      I2 => blk00000001_sig00000205,
      I3 => blk00000001_sig00000225,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000492
    );
  blk00000001_blk0000026a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000244,
      I1 => blk00000001_sig000001e4,
      I2 => blk00000001_sig00000204,
      I3 => blk00000001_sig00000224,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000491
    );
  blk00000001_blk00000269 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000243,
      I1 => blk00000001_sig000001e3,
      I2 => blk00000001_sig00000203,
      I3 => blk00000001_sig00000223,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000490
    );
  blk00000001_blk00000268 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000242,
      I1 => blk00000001_sig000001e2,
      I2 => blk00000001_sig00000202,
      I3 => blk00000001_sig00000222,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048f
    );
  blk00000001_blk00000267 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000241,
      I1 => blk00000001_sig000001e1,
      I2 => blk00000001_sig00000201,
      I3 => blk00000001_sig00000221,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048e
    );
  blk00000001_blk00000266 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048d,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000407
    );
  blk00000001_blk00000265 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048c,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000406
    );
  blk00000001_blk00000264 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048b,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000405
    );
  blk00000001_blk00000263 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000048a,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000404
    );
  blk00000001_blk00000262 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000489,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000403
    );
  blk00000001_blk00000261 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000488,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000402
    );
  blk00000001_blk00000260 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000487,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000401
    );
  blk00000001_blk0000025f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000486,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000400
    );
  blk00000001_blk0000025e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000485,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003ff
    );
  blk00000001_blk0000025d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000484,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003fe
    );
  blk00000001_blk0000025c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000483,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003fd
    );
  blk00000001_blk0000025b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000482,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003fc
    );
  blk00000001_blk0000025a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000481,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003fb
    );
  blk00000001_blk00000259 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000480,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003fa
    );
  blk00000001_blk00000258 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f9
    );
  blk00000001_blk00000257 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000003f8
    );
  blk00000001_blk00000256 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000200,
      I1 => blk00000001_sig00000220,
      I2 => blk00000001_sig00000240,
      I3 => blk00000001_sig00000260,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048d
    );
  blk00000001_blk00000255 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001ff,
      I1 => blk00000001_sig0000021f,
      I2 => blk00000001_sig0000023f,
      I3 => blk00000001_sig0000025f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048c
    );
  blk00000001_blk00000254 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fe,
      I1 => blk00000001_sig0000021e,
      I2 => blk00000001_sig0000023e,
      I3 => blk00000001_sig0000025e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048b
    );
  blk00000001_blk00000253 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fd,
      I1 => blk00000001_sig0000021d,
      I2 => blk00000001_sig0000023d,
      I3 => blk00000001_sig0000025d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000048a
    );
  blk00000001_blk00000252 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fc,
      I1 => blk00000001_sig0000021c,
      I2 => blk00000001_sig0000023c,
      I3 => blk00000001_sig0000025c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000489
    );
  blk00000001_blk00000251 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fb,
      I1 => blk00000001_sig0000021b,
      I2 => blk00000001_sig0000023b,
      I3 => blk00000001_sig0000025b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000488
    );
  blk00000001_blk00000250 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001fa,
      I1 => blk00000001_sig0000021a,
      I2 => blk00000001_sig0000023a,
      I3 => blk00000001_sig0000025a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000487
    );
  blk00000001_blk0000024f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f9,
      I1 => blk00000001_sig00000219,
      I2 => blk00000001_sig00000239,
      I3 => blk00000001_sig00000259,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000486
    );
  blk00000001_blk0000024e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f8,
      I1 => blk00000001_sig00000218,
      I2 => blk00000001_sig00000238,
      I3 => blk00000001_sig00000258,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000485
    );
  blk00000001_blk0000024d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f7,
      I1 => blk00000001_sig00000217,
      I2 => blk00000001_sig00000237,
      I3 => blk00000001_sig00000257,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000484
    );
  blk00000001_blk0000024c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f6,
      I1 => blk00000001_sig00000216,
      I2 => blk00000001_sig00000236,
      I3 => blk00000001_sig00000256,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000483
    );
  blk00000001_blk0000024b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f5,
      I1 => blk00000001_sig00000215,
      I2 => blk00000001_sig00000235,
      I3 => blk00000001_sig00000255,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000482
    );
  blk00000001_blk0000024a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f4,
      I1 => blk00000001_sig00000214,
      I2 => blk00000001_sig00000234,
      I3 => blk00000001_sig00000254,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000481
    );
  blk00000001_blk00000249 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f3,
      I1 => blk00000001_sig00000213,
      I2 => blk00000001_sig00000233,
      I3 => blk00000001_sig00000253,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000480
    );
  blk00000001_blk00000248 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f2,
      I1 => blk00000001_sig00000212,
      I2 => blk00000001_sig00000232,
      I3 => blk00000001_sig00000252,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047f
    );
  blk00000001_blk00000247 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig000001f1,
      I1 => blk00000001_sig00000211,
      I2 => blk00000001_sig00000231,
      I3 => blk00000001_sig00000251,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047e
    );
  blk00000001_blk00000246 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047d,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e7
    );
  blk00000001_blk00000245 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047c,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e6
    );
  blk00000001_blk00000244 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047b,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e5
    );
  blk00000001_blk00000243 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000047a,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e4
    );
  blk00000001_blk00000242 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000479,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e3
    );
  blk00000001_blk00000241 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000478,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e2
    );
  blk00000001_blk00000240 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000477,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e1
    );
  blk00000001_blk0000023f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000476,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007e0
    );
  blk00000001_blk0000023e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000475,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007df
    );
  blk00000001_blk0000023d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000474,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007de
    );
  blk00000001_blk0000023c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000473,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007dd
    );
  blk00000001_blk0000023b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000472,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007dc
    );
  blk00000001_blk0000023a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000471,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007db
    );
  blk00000001_blk00000239 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000470,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007da
    );
  blk00000001_blk00000238 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d9
    );
  blk00000001_blk00000237 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000007d8
    );
  blk00000001_blk00000236 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000220,
      I1 => blk00000001_sig00000240,
      I2 => blk00000001_sig00000260,
      I3 => blk00000001_sig00000200,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047d
    );
  blk00000001_blk00000235 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021f,
      I1 => blk00000001_sig0000023f,
      I2 => blk00000001_sig0000025f,
      I3 => blk00000001_sig000001ff,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047c
    );
  blk00000001_blk00000234 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021e,
      I1 => blk00000001_sig0000023e,
      I2 => blk00000001_sig0000025e,
      I3 => blk00000001_sig000001fe,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047b
    );
  blk00000001_blk00000233 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021d,
      I1 => blk00000001_sig0000023d,
      I2 => blk00000001_sig0000025d,
      I3 => blk00000001_sig000001fd,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000047a
    );
  blk00000001_blk00000232 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021c,
      I1 => blk00000001_sig0000023c,
      I2 => blk00000001_sig0000025c,
      I3 => blk00000001_sig000001fc,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000479
    );
  blk00000001_blk00000231 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021b,
      I1 => blk00000001_sig0000023b,
      I2 => blk00000001_sig0000025b,
      I3 => blk00000001_sig000001fb,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000478
    );
  blk00000001_blk00000230 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000021a,
      I1 => blk00000001_sig0000023a,
      I2 => blk00000001_sig0000025a,
      I3 => blk00000001_sig000001fa,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000477
    );
  blk00000001_blk0000022f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000219,
      I1 => blk00000001_sig00000239,
      I2 => blk00000001_sig00000259,
      I3 => blk00000001_sig000001f9,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000476
    );
  blk00000001_blk0000022e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000218,
      I1 => blk00000001_sig00000238,
      I2 => blk00000001_sig00000258,
      I3 => blk00000001_sig000001f8,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000475
    );
  blk00000001_blk0000022d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000217,
      I1 => blk00000001_sig00000237,
      I2 => blk00000001_sig00000257,
      I3 => blk00000001_sig000001f7,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000474
    );
  blk00000001_blk0000022c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000216,
      I1 => blk00000001_sig00000236,
      I2 => blk00000001_sig00000256,
      I3 => blk00000001_sig000001f6,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000473
    );
  blk00000001_blk0000022b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000215,
      I1 => blk00000001_sig00000235,
      I2 => blk00000001_sig00000255,
      I3 => blk00000001_sig000001f5,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000472
    );
  blk00000001_blk0000022a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000214,
      I1 => blk00000001_sig00000234,
      I2 => blk00000001_sig00000254,
      I3 => blk00000001_sig000001f4,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000471
    );
  blk00000001_blk00000229 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000213,
      I1 => blk00000001_sig00000233,
      I2 => blk00000001_sig00000253,
      I3 => blk00000001_sig000001f3,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000470
    );
  blk00000001_blk00000228 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000212,
      I1 => blk00000001_sig00000232,
      I2 => blk00000001_sig00000252,
      I3 => blk00000001_sig000001f2,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046f
    );
  blk00000001_blk00000227 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000211,
      I1 => blk00000001_sig00000231,
      I2 => blk00000001_sig00000251,
      I3 => blk00000001_sig000001f1,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046e
    );
  blk00000001_blk00000226 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046d,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000085a
    );
  blk00000001_blk00000225 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046c,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000859
    );
  blk00000001_blk00000224 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046b,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000858
    );
  blk00000001_blk00000223 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000046a,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000857
    );
  blk00000001_blk00000222 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000469,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000856
    );
  blk00000001_blk00000221 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000468,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000855
    );
  blk00000001_blk00000220 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000467,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000854
    );
  blk00000001_blk0000021f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000466,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000853
    );
  blk00000001_blk0000021e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000465,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000852
    );
  blk00000001_blk0000021d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000464,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000851
    );
  blk00000001_blk0000021c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000463,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig00000850
    );
  blk00000001_blk0000021b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000462,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084f
    );
  blk00000001_blk0000021a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000461,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084e
    );
  blk00000001_blk00000219 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000460,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084d
    );
  blk00000001_blk00000218 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084c
    );
  blk00000001_blk00000217 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig0000084b
    );
  blk00000001_blk00000216 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000240,
      I1 => blk00000001_sig00000260,
      I2 => blk00000001_sig00000200,
      I3 => blk00000001_sig00000220,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046d
    );
  blk00000001_blk00000215 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023f,
      I1 => blk00000001_sig0000025f,
      I2 => blk00000001_sig000001ff,
      I3 => blk00000001_sig0000021f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046c
    );
  blk00000001_blk00000214 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023e,
      I1 => blk00000001_sig0000025e,
      I2 => blk00000001_sig000001fe,
      I3 => blk00000001_sig0000021e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046b
    );
  blk00000001_blk00000213 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023d,
      I1 => blk00000001_sig0000025d,
      I2 => blk00000001_sig000001fd,
      I3 => blk00000001_sig0000021d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000046a
    );
  blk00000001_blk00000212 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023c,
      I1 => blk00000001_sig0000025c,
      I2 => blk00000001_sig000001fc,
      I3 => blk00000001_sig0000021c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000469
    );
  blk00000001_blk00000211 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023b,
      I1 => blk00000001_sig0000025b,
      I2 => blk00000001_sig000001fb,
      I3 => blk00000001_sig0000021b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000468
    );
  blk00000001_blk00000210 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000023a,
      I1 => blk00000001_sig0000025a,
      I2 => blk00000001_sig000001fa,
      I3 => blk00000001_sig0000021a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000467
    );
  blk00000001_blk0000020f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000239,
      I1 => blk00000001_sig00000259,
      I2 => blk00000001_sig000001f9,
      I3 => blk00000001_sig00000219,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000466
    );
  blk00000001_blk0000020e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000238,
      I1 => blk00000001_sig00000258,
      I2 => blk00000001_sig000001f8,
      I3 => blk00000001_sig00000218,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000465
    );
  blk00000001_blk0000020d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000237,
      I1 => blk00000001_sig00000257,
      I2 => blk00000001_sig000001f7,
      I3 => blk00000001_sig00000217,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000464
    );
  blk00000001_blk0000020c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000236,
      I1 => blk00000001_sig00000256,
      I2 => blk00000001_sig000001f6,
      I3 => blk00000001_sig00000216,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000463
    );
  blk00000001_blk0000020b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000235,
      I1 => blk00000001_sig00000255,
      I2 => blk00000001_sig000001f5,
      I3 => blk00000001_sig00000215,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000462
    );
  blk00000001_blk0000020a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000234,
      I1 => blk00000001_sig00000254,
      I2 => blk00000001_sig000001f4,
      I3 => blk00000001_sig00000214,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000461
    );
  blk00000001_blk00000209 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000233,
      I1 => blk00000001_sig00000253,
      I2 => blk00000001_sig000001f3,
      I3 => blk00000001_sig00000213,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000460
    );
  blk00000001_blk00000208 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000232,
      I1 => blk00000001_sig00000252,
      I2 => blk00000001_sig000001f2,
      I3 => blk00000001_sig00000212,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045f
    );
  blk00000001_blk00000207 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000231,
      I1 => blk00000001_sig00000251,
      I2 => blk00000001_sig000001f1,
      I3 => blk00000001_sig00000211,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045e
    );
  blk00000001_blk00000206 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045d,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008cf
    );
  blk00000001_blk00000205 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045c,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008ce
    );
  blk00000001_blk00000204 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045b,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008cd
    );
  blk00000001_blk00000203 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000045a,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008cc
    );
  blk00000001_blk00000202 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000459,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008cb
    );
  blk00000001_blk00000201 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000458,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008ca
    );
  blk00000001_blk00000200 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000457,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c9
    );
  blk00000001_blk000001ff : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000456,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c8
    );
  blk00000001_blk000001fe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000455,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c7
    );
  blk00000001_blk000001fd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000454,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c6
    );
  blk00000001_blk000001fc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000453,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c5
    );
  blk00000001_blk000001fb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000452,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c4
    );
  blk00000001_blk000001fa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000451,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c3
    );
  blk00000001_blk000001f9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig00000450,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c2
    );
  blk00000001_blk000001f8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000044f,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c1
    );
  blk00000001_blk000001f7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001ae,
      D => blk00000001_sig0000044e,
      R => blk00000001_sig000001a4,
      Q => blk00000001_sig000008c0
    );
  blk00000001_blk000001f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000260,
      I1 => blk00000001_sig00000200,
      I2 => blk00000001_sig00000220,
      I3 => blk00000001_sig00000240,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045d
    );
  blk00000001_blk000001f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025f,
      I1 => blk00000001_sig000001ff,
      I2 => blk00000001_sig0000021f,
      I3 => blk00000001_sig0000023f,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045c
    );
  blk00000001_blk000001f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025e,
      I1 => blk00000001_sig000001fe,
      I2 => blk00000001_sig0000021e,
      I3 => blk00000001_sig0000023e,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045b
    );
  blk00000001_blk000001f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025d,
      I1 => blk00000001_sig000001fd,
      I2 => blk00000001_sig0000021d,
      I3 => blk00000001_sig0000023d,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000045a
    );
  blk00000001_blk000001f2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025c,
      I1 => blk00000001_sig000001fc,
      I2 => blk00000001_sig0000021c,
      I3 => blk00000001_sig0000023c,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000459
    );
  blk00000001_blk000001f1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025b,
      I1 => blk00000001_sig000001fb,
      I2 => blk00000001_sig0000021b,
      I3 => blk00000001_sig0000023b,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000458
    );
  blk00000001_blk000001f0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig0000025a,
      I1 => blk00000001_sig000001fa,
      I2 => blk00000001_sig0000021a,
      I3 => blk00000001_sig0000023a,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000457
    );
  blk00000001_blk000001ef : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000259,
      I1 => blk00000001_sig000001f9,
      I2 => blk00000001_sig00000219,
      I3 => blk00000001_sig00000239,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000456
    );
  blk00000001_blk000001ee : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000258,
      I1 => blk00000001_sig000001f8,
      I2 => blk00000001_sig00000218,
      I3 => blk00000001_sig00000238,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000455
    );
  blk00000001_blk000001ed : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000257,
      I1 => blk00000001_sig000001f7,
      I2 => blk00000001_sig00000217,
      I3 => blk00000001_sig00000237,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000454
    );
  blk00000001_blk000001ec : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000256,
      I1 => blk00000001_sig000001f6,
      I2 => blk00000001_sig00000216,
      I3 => blk00000001_sig00000236,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000453
    );
  blk00000001_blk000001eb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000255,
      I1 => blk00000001_sig000001f5,
      I2 => blk00000001_sig00000215,
      I3 => blk00000001_sig00000235,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000452
    );
  blk00000001_blk000001ea : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000254,
      I1 => blk00000001_sig000001f4,
      I2 => blk00000001_sig00000214,
      I3 => blk00000001_sig00000234,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000451
    );
  blk00000001_blk000001e9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000253,
      I1 => blk00000001_sig000001f3,
      I2 => blk00000001_sig00000213,
      I3 => blk00000001_sig00000233,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig00000450
    );
  blk00000001_blk000001e8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000252,
      I1 => blk00000001_sig000001f2,
      I2 => blk00000001_sig00000212,
      I3 => blk00000001_sig00000232,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000044f
    );
  blk00000001_blk000001e7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_sig00000251,
      I1 => blk00000001_sig000001f1,
      I2 => blk00000001_sig00000211,
      I3 => blk00000001_sig00000231,
      I4 => blk00000001_sig000001b7,
      I5 => blk00000001_sig000001b8,
      O => blk00000001_sig0000044e
    );
  blk00000001_blk000001e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000044d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041e
    );
  blk00000001_blk000001e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000044c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041f
    );
  blk00000001_blk000001e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000044b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000420
    );
  blk00000001_blk000001e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000044a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000421
    );
  blk00000001_blk000001e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000449,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000422
    );
  blk00000001_blk000001e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000448,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000423
    );
  blk00000001_blk000001e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000447,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000424
    );
  blk00000001_blk000001df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000446,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000425
    );
  blk00000001_blk000001de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000445,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000426
    );
  blk00000001_blk000001dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000444,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000427
    );
  blk00000001_blk000001dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000443,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000428
    );
  blk00000001_blk000001db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000442,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000429
    );
  blk00000001_blk000001da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000441,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000042a
    );
  blk00000001_blk000001d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000440,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000042b
    );
  blk00000001_blk000001d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000042c
    );
  blk00000001_blk000001d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000042d
    );
  blk00000001_blk000001d6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000067,
      Q => blk00000001_sig0000044d
    );
  blk00000001_blk000001d5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000066,
      Q => blk00000001_sig0000044c
    );
  blk00000001_blk000001d4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000065,
      Q => blk00000001_sig0000044b
    );
  blk00000001_blk000001d3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000064,
      Q => blk00000001_sig0000044a
    );
  blk00000001_blk000001d2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000063,
      Q => blk00000001_sig00000449
    );
  blk00000001_blk000001d1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000062,
      Q => blk00000001_sig00000448
    );
  blk00000001_blk000001d0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000061,
      Q => blk00000001_sig00000447
    );
  blk00000001_blk000001cf : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000060,
      Q => blk00000001_sig00000446
    );
  blk00000001_blk000001ce : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005f,
      Q => blk00000001_sig00000445
    );
  blk00000001_blk000001cd : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005e,
      Q => blk00000001_sig00000444
    );
  blk00000001_blk000001cc : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005d,
      Q => blk00000001_sig00000443
    );
  blk00000001_blk000001cb : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005c,
      Q => blk00000001_sig00000442
    );
  blk00000001_blk000001ca : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005b,
      Q => blk00000001_sig00000441
    );
  blk00000001_blk000001c9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000005a,
      Q => blk00000001_sig00000440
    );
  blk00000001_blk000001c8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000059,
      Q => blk00000001_sig0000043f
    );
  blk00000001_blk000001c7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000058,
      Q => blk00000001_sig0000043e
    );
  blk00000001_blk000001c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043d,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000040e
    );
  blk00000001_blk000001c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043c,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000040f
    );
  blk00000001_blk000001c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043b,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000410
    );
  blk00000001_blk000001c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000043a,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000411
    );
  blk00000001_blk000001c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000439,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000412
    );
  blk00000001_blk000001c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000438,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000413
    );
  blk00000001_blk000001c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000437,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000414
    );
  blk00000001_blk000001bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000436,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000415
    );
  blk00000001_blk000001be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000435,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000416
    );
  blk00000001_blk000001bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000434,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000417
    );
  blk00000001_blk000001bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000433,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000418
    );
  blk00000001_blk000001bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000432,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig00000419
    );
  blk00000001_blk000001ba : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000431,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041a
    );
  blk00000001_blk000001b9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000430,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041b
    );
  blk00000001_blk000001b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000042f,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041c
    );
  blk00000001_blk000001b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000042e,
      R => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      Q => blk00000001_sig0000041d
    );
  blk00000001_blk000001b6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000077,
      Q => blk00000001_sig0000043d
    );
  blk00000001_blk000001b5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000076,
      Q => blk00000001_sig0000043c
    );
  blk00000001_blk000001b4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000075,
      Q => blk00000001_sig0000043b
    );
  blk00000001_blk000001b3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000074,
      Q => blk00000001_sig0000043a
    );
  blk00000001_blk000001b2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000073,
      Q => blk00000001_sig00000439
    );
  blk00000001_blk000001b1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000072,
      Q => blk00000001_sig00000438
    );
  blk00000001_blk000001b0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000071,
      Q => blk00000001_sig00000437
    );
  blk00000001_blk000001af : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000070,
      Q => blk00000001_sig00000436
    );
  blk00000001_blk000001ae : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006f,
      Q => blk00000001_sig00000435
    );
  blk00000001_blk000001ad : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006e,
      Q => blk00000001_sig00000434
    );
  blk00000001_blk000001ac : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006d,
      Q => blk00000001_sig00000433
    );
  blk00000001_blk000001ab : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006c,
      Q => blk00000001_sig00000432
    );
  blk00000001_blk000001aa : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006b,
      Q => blk00000001_sig00000431
    );
  blk00000001_blk000001a9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig0000006a,
      Q => blk00000001_sig00000430
    );
  blk00000001_blk000001a8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000069,
      Q => blk00000001_sig0000042f
    );
  blk00000001_blk000001a7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_sig000000c0,
      A1 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A2 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      A3 => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000068,
      Q => blk00000001_sig0000042e
    );
  blk00000001_blk000001a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig0000007d,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig00000408
    );
  blk00000001_blk000001a5 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig0000007c,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig00000409
    );
  blk00000001_blk000001a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig0000007b,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig0000040a
    );
  blk00000001_blk000001a3 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig0000007a,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig0000040b
    );
  blk00000001_blk000001a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig00000079,
      R => blk00000001_sig0000008d,
      Q => blk00000001_sig0000040c
    );
  blk00000001_blk000001a1 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig00000078,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig0000040d
    );
  blk00000001_blk000001a0 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000002e3,
      D => blk00000001_sig0000008c,
      S => blk00000001_sig0000008d,
      Q => blk00000001_sig000002e4
    );
  blk00000001_blk0000019f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig000002e4,
      Q => blk00000001_sig000001e0
    );
  blk00000001_blk0000019e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig00000408,
      Q => blk00000001_sig000001da
    );
  blk00000001_blk0000019d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig00000409,
      Q => blk00000001_sig000001db
    );
  blk00000001_blk0000019c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig0000040a,
      Q => blk00000001_sig000001dc
    );
  blk00000001_blk0000019b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig0000040b,
      Q => blk00000001_sig000001dd
    );
  blk00000001_blk0000019a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig0000040c,
      Q => blk00000001_sig000001de
    );
  blk00000001_blk00000199 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000001a5,
      D => blk00000001_sig0000040d,
      Q => blk00000001_sig000001df
    );
  blk00000001_blk000000b0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tlast,
      Q => blk00000001_sig00000183
    );
  blk00000001_blk000000af : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(0),
      Q => blk00000001_sig00000184
    );
  blk00000001_blk000000ae : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(1),
      Q => blk00000001_sig00000185
    );
  blk00000001_blk000000ad : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(2),
      Q => blk00000001_sig00000186
    );
  blk00000001_blk000000ac : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(3),
      Q => blk00000001_sig00000187
    );
  blk00000001_blk000000ab : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(4),
      Q => blk00000001_sig00000188
    );
  blk00000001_blk000000aa : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(5),
      Q => blk00000001_sig00000189
    );
  blk00000001_blk000000a9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(6),
      Q => blk00000001_sig0000018a
    );
  blk00000001_blk000000a8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(7),
      Q => blk00000001_sig0000018b
    );
  blk00000001_blk000000a7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(8),
      Q => blk00000001_sig0000018c
    );
  blk00000001_blk000000a6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(9),
      Q => blk00000001_sig0000018d
    );
  blk00000001_blk000000a5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(10),
      Q => blk00000001_sig0000018e
    );
  blk00000001_blk000000a4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(11),
      Q => blk00000001_sig0000018f
    );
  blk00000001_blk000000a3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(12),
      Q => blk00000001_sig00000190
    );
  blk00000001_blk000000a2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(13),
      Q => blk00000001_sig00000191
    );
  blk00000001_blk000000a1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(14),
      Q => blk00000001_sig00000192
    );
  blk00000001_blk000000a0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(15),
      Q => blk00000001_sig00000193
    );
  blk00000001_blk0000009f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(16),
      Q => blk00000001_sig00000194
    );
  blk00000001_blk0000009e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(17),
      Q => blk00000001_sig00000195
    );
  blk00000001_blk0000009d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(18),
      Q => blk00000001_sig00000196
    );
  blk00000001_blk0000009c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(19),
      Q => blk00000001_sig00000197
    );
  blk00000001_blk0000009b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(20),
      Q => blk00000001_sig00000198
    );
  blk00000001_blk0000009a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(21),
      Q => blk00000001_sig00000199
    );
  blk00000001_blk00000099 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(22),
      Q => blk00000001_sig0000019a
    );
  blk00000001_blk00000098 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(23),
      Q => blk00000001_sig0000019b
    );
  blk00000001_blk00000097 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(24),
      Q => blk00000001_sig0000019c
    );
  blk00000001_blk00000096 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(25),
      Q => blk00000001_sig0000019d
    );
  blk00000001_blk00000095 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(26),
      Q => blk00000001_sig0000019e
    );
  blk00000001_blk00000094 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(27),
      Q => blk00000001_sig0000019f
    );
  blk00000001_blk00000093 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(28),
      Q => blk00000001_sig000001a0
    );
  blk00000001_blk00000092 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(29),
      Q => blk00000001_sig000001a1
    );
  blk00000001_blk00000091 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(30),
      Q => blk00000001_sig000001a2
    );
  blk00000001_blk00000090 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(31),
      Q => blk00000001_sig000001a3
    );
  blk00000001_blk0000008f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig0000017f,
      Q => NlwRenamedSig_OI_s_axis_data_tready
    );
  blk00000001_blk0000008e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000180,
      Q => blk00000001_sig00000181
    );
  blk00000001_blk0000008d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000faa,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013b
    );
  blk00000001_blk0000008c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fab,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013c
    );
  blk00000001_blk0000008b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fac,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013d
    );
  blk00000001_blk0000008a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fad,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013e
    );
  blk00000001_blk00000089 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fae,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000013f
    );
  blk00000001_blk00000088 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000faf,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000140
    );
  blk00000001_blk00000087 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb0,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000141
    );
  blk00000001_blk00000086 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb1,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000142
    );
  blk00000001_blk00000085 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb2,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000143
    );
  blk00000001_blk00000084 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb3,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000144
    );
  blk00000001_blk00000083 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb4,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000145
    );
  blk00000001_blk00000082 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb5,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000146
    );
  blk00000001_blk00000081 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb6,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000147
    );
  blk00000001_blk00000080 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb7,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000148
    );
  blk00000001_blk0000007f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb8,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000149
    );
  blk00000001_blk0000007e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fb9,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014a
    );
  blk00000001_blk0000007d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fba,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014b
    );
  blk00000001_blk0000007c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fbb,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014c
    );
  blk00000001_blk0000007b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fbc,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014d
    );
  blk00000001_blk0000007a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fbd,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014e
    );
  blk00000001_blk00000079 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fbe,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000014f
    );
  blk00000001_blk00000078 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fbf,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000150
    );
  blk00000001_blk00000077 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc0,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000151
    );
  blk00000001_blk00000076 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc1,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000152
    );
  blk00000001_blk00000075 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc2,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000153
    );
  blk00000001_blk00000074 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc3,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000154
    );
  blk00000001_blk00000073 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc4,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000155
    );
  blk00000001_blk00000072 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc5,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000156
    );
  blk00000001_blk00000071 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc6,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000157
    );
  blk00000001_blk00000070 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc7,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000158
    );
  blk00000001_blk0000006f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc8,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000159
    );
  blk00000001_blk0000006e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fc9,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000015a
    );
  blk00000001_blk0000006d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000fa9,
      D => blk00000001_sig00000fca,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000015b
    );
  blk00000001_blk0000006c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000118,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000102
    );
  blk00000001_blk0000006b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000119,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000067
    );
  blk00000001_blk0000006a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011a,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000066
    );
  blk00000001_blk00000069 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011b,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000065
    );
  blk00000001_blk00000068 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011c,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000064
    );
  blk00000001_blk00000067 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011d,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000063
    );
  blk00000001_blk00000066 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011e,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000062
    );
  blk00000001_blk00000065 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000011f,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000061
    );
  blk00000001_blk00000064 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000120,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000060
    );
  blk00000001_blk00000063 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000121,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005f
    );
  blk00000001_blk00000062 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000122,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005e
    );
  blk00000001_blk00000061 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000123,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005d
    );
  blk00000001_blk00000060 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000124,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005c
    );
  blk00000001_blk0000005f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000125,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005b
    );
  blk00000001_blk0000005e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000126,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000005a
    );
  blk00000001_blk0000005d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000127,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000059
    );
  blk00000001_blk0000005c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000128,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000058
    );
  blk00000001_blk0000005b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000129,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000077
    );
  blk00000001_blk0000005a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012a,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000076
    );
  blk00000001_blk00000059 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012b,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000075
    );
  blk00000001_blk00000058 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012c,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000074
    );
  blk00000001_blk00000057 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012d,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000073
    );
  blk00000001_blk00000056 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012e,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000072
    );
  blk00000001_blk00000055 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig0000012f,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000071
    );
  blk00000001_blk00000054 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000130,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000070
    );
  blk00000001_blk00000053 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000131,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006f
    );
  blk00000001_blk00000052 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000132,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006e
    );
  blk00000001_blk00000051 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000133,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006d
    );
  blk00000001_blk00000050 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000134,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006c
    );
  blk00000001_blk0000004f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000135,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006b
    );
  blk00000001_blk0000004e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000136,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000006a
    );
  blk00000001_blk0000004d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000137,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000069
    );
  blk00000001_blk0000004c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000116,
      D => blk00000001_sig00000138,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000068
    );
  blk00000001_blk00000024 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(0),
      Q => blk00000001_sig0000010f
    );
  blk00000001_blk00000023 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(1),
      Q => blk00000001_sig00000110
    );
  blk00000001_blk00000022 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(2),
      Q => blk00000001_sig00000111
    );
  blk00000001_blk00000021 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(3),
      Q => blk00000001_sig00000112
    );
  blk00000001_blk00000020 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(4),
      Q => blk00000001_sig00000113
    );
  blk00000001_blk0000001f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(5),
      Q => blk00000001_sig00000114
    );
  blk00000001_blk0000001e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(6),
      Q => blk00000001_sig00000115
    );
  blk00000001_blk0000001d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig0000010b,
      Q => NlwRenamedSig_OI_s_axis_config_tready
    );
  blk00000001_blk0000001c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig0000010c,
      Q => blk00000001_sig0000010d
    );
  blk00000001_blk0000001b : FDR
    port map (
      C => aclk,
      D => blk00000001_sig000000cf,
      R => blk00000001_sig000000cc,
      Q => blk00000001_sig0000008e
    );
  blk00000001_blk0000001a : FDS
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig000000cc,
      Q => blk00000001_sig000000f9
    );
  blk00000001_blk00000019 : FDS
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000f9,
      S => blk00000001_sig000000cc,
      Q => blk00000001_sig000000f8
    );
  blk00000001_blk00000018 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000cd,
      R => blk00000001_sig000000f8,
      Q => event_tlast_unexpected
    );
  blk00000001_blk00000017 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000d2,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000fa
    );
  blk00000001_blk00000016 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000d1,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000008b
    );
  blk00000001_blk00000015 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000be,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f4
    );
  blk00000001_blk00000014 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000d3,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig0000008d
    );
  blk00000001_blk00000013 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000d0,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e2
    );
  blk00000001_blk00000012 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig0000008a,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e1
    );
  blk00000001_blk00000011 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000d5,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000df
    );
  blk00000001_blk00000010 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000ce,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e0
    );
  blk00000001_blk0000000f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000d4,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000de
    );
  blk00000001_blk0000000e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig000000dd,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e3
    );
  blk00000001_blk0000000d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_sig00000103,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000f5
    );
  blk00000001_blk0000000c : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000104,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e4
    );
  blk00000001_blk0000000b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000105,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e5
    );
  blk00000001_blk0000000a : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000106,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e6
    );
  blk00000001_blk00000009 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000107,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e7
    );
  blk00000001_blk00000008 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000108,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e8
    );
  blk00000001_blk00000007 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig00000109,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000e9
    );
  blk00000001_blk00000006 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig000000f7,
      D => blk00000001_sig0000010a,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig000000ea
    );
  blk00000001_blk00000005 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000c8,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000fb
    );
  blk00000001_blk00000004 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000c7,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig000000fc
    );
  blk00000001_blk00000003 : GND
    port map (
      G => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000002 : VCC
    port map (
      P => blk00000001_sig000000c0
    );
  blk00000001_blk00000025_blk0000004b : INV
    port map (
      I => blk00000001_blk00000025_sig00000fe9,
      O => blk00000001_blk00000025_sig00000ff6
    );
  blk00000001_blk00000025_blk0000004a : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000fe9,
      I1 => blk00000001_sig000000f7,
      O => blk00000001_blk00000025_sig00001004
    );
  blk00000001_blk00000025_blk00000049 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000fea,
      I1 => blk00000001_blk00000025_sig00000fe9,
      I2 => blk00000001_sig000000f7,
      O => blk00000001_blk00000025_sig00001002
    );
  blk00000001_blk00000025_blk00000048 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000feb,
      I1 => blk00000001_blk00000025_sig00000fe9,
      I2 => blk00000001_sig000000f7,
      O => blk00000001_blk00000025_sig00001000
    );
  blk00000001_blk00000025_blk00000047 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000fec,
      I1 => blk00000001_blk00000025_sig00000fe9,
      I2 => blk00000001_sig000000f7,
      O => blk00000001_blk00000025_sig00000ffe
    );
  blk00000001_blk00000025_blk00000046 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000fed,
      I1 => blk00000001_blk00000025_sig00000fe9,
      I2 => blk00000001_sig000000f7,
      O => blk00000001_blk00000025_sig00000ffc
    );
  blk00000001_blk00000025_blk00000045 : LUT6
    generic map(
      INIT => X"8AAA8A8AAABAAAAA"
    )
    port map (
      I0 => blk00000001_sig0000010e,
      I1 => blk00000001_blk00000025_sig00001005,
      I2 => blk00000001_blk00000025_sig00000fea,
      I3 => blk00000001_blk00000025_sig00000fe9,
      I4 => blk00000001_sig000000f7,
      I5 => blk00000001_sig0000010d,
      O => blk00000001_blk00000025_sig00000ff5
    );
  blk00000001_blk00000025_blk00000044 : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_blk00000025_sig00000fed,
      I1 => blk00000001_blk00000025_sig00000feb,
      I2 => blk00000001_blk00000025_sig00000fec,
      O => blk00000001_blk00000025_sig00001005
    );
  blk00000001_blk00000025_blk00000043 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000115,
      Q => blk00000001_blk00000025_sig00000fee,
      Q15 => NLW_blk00000001_blk00000025_blk00000043_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000042 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000114,
      Q => blk00000001_blk00000025_sig00000fef,
      Q15 => NLW_blk00000001_blk00000025_blk00000042_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000041 : XORCY
    port map (
      CI => blk00000001_blk00000025_sig00001003,
      LI => blk00000001_blk00000025_sig00001004,
      O => blk00000001_blk00000025_sig00000ffb
    );
  blk00000001_blk00000025_blk00000040 : XORCY
    port map (
      CI => blk00000001_blk00000025_sig00001001,
      LI => blk00000001_blk00000025_sig00001002,
      O => blk00000001_blk00000025_sig00000ffa
    );
  blk00000001_blk00000025_blk0000003f : MUXCY
    port map (
      CI => blk00000001_blk00000025_sig00001001,
      DI => blk00000001_blk00000025_sig00000fea,
      S => blk00000001_blk00000025_sig00001002,
      O => blk00000001_blk00000025_sig00001003
    );
  blk00000001_blk00000025_blk0000003e : XORCY
    port map (
      CI => blk00000001_blk00000025_sig00000fff,
      LI => blk00000001_blk00000025_sig00001000,
      O => blk00000001_blk00000025_sig00000ff9
    );
  blk00000001_blk00000025_blk0000003d : MUXCY
    port map (
      CI => blk00000001_blk00000025_sig00000fff,
      DI => blk00000001_blk00000025_sig00000feb,
      S => blk00000001_blk00000025_sig00001000,
      O => blk00000001_blk00000025_sig00001001
    );
  blk00000001_blk00000025_blk0000003c : XORCY
    port map (
      CI => blk00000001_blk00000025_sig00000ffd,
      LI => blk00000001_blk00000025_sig00000ffe,
      O => blk00000001_blk00000025_sig00000ff8
    );
  blk00000001_blk00000025_blk0000003b : MUXCY
    port map (
      CI => blk00000001_blk00000025_sig00000ffd,
      DI => blk00000001_blk00000025_sig00000fec,
      S => blk00000001_blk00000025_sig00000ffe,
      O => blk00000001_blk00000025_sig00000fff
    );
  blk00000001_blk00000025_blk0000003a : XORCY
    port map (
      CI => blk00000001_sig0000010d,
      LI => blk00000001_blk00000025_sig00000ffc,
      O => blk00000001_blk00000025_sig00000ff7
    );
  blk00000001_blk00000025_blk00000039 : MUXCY
    port map (
      CI => blk00000001_sig0000010d,
      DI => blk00000001_blk00000025_sig00000fed,
      S => blk00000001_blk00000025_sig00000ffc,
      O => blk00000001_blk00000025_sig00000ffd
    );
  blk00000001_blk00000025_blk00000038 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000112,
      Q => blk00000001_blk00000025_sig00000ff1,
      Q15 => NLW_blk00000001_blk00000025_blk00000038_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000037 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000111,
      Q => blk00000001_blk00000025_sig00000ff2,
      Q15 => NLW_blk00000001_blk00000025_blk00000037_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000036 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000113,
      Q => blk00000001_blk00000025_sig00000ff0,
      Q15 => NLW_blk00000001_blk00000025_blk00000036_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000035 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig0000010f,
      Q => blk00000001_blk00000025_sig00000ff4,
      Q15 => NLW_blk00000001_blk00000025_blk00000035_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000034 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000025_sig00000fed,
      A1 => blk00000001_blk00000025_sig00000fec,
      A2 => blk00000001_blk00000025_sig00000feb,
      A3 => blk00000001_blk00000025_sig00000fea,
      CE => blk00000001_sig0000010d,
      CLK => aclk,
      D => blk00000001_sig00000110,
      Q => blk00000001_blk00000025_sig00000ff3,
      Q15 => NLW_blk00000001_blk00000025_blk00000034_Q15_UNCONNECTED
    );
  blk00000001_blk00000025_blk00000033 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ffb,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk00000025_sig00000fe9
    );
  blk00000001_blk00000025_blk00000032 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ffa,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk00000025_sig00000fea
    );
  blk00000001_blk00000025_blk00000031 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff9,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk00000025_sig00000feb
    );
  blk00000001_blk00000025_blk00000030 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff8,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk00000025_sig00000fec
    );
  blk00000001_blk00000025_blk0000002f : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff7,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk00000025_sig00000fed
    );
  blk00000001_blk00000025_blk0000002e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000fee,
      Q => blk00000001_sig0000010a
    );
  blk00000001_blk00000025_blk0000002d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000fef,
      Q => blk00000001_sig00000109
    );
  blk00000001_blk00000025_blk0000002c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff0,
      Q => blk00000001_sig00000108
    );
  blk00000001_blk00000025_blk0000002b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff1,
      Q => blk00000001_sig00000107
    );
  blk00000001_blk00000025_blk0000002a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff2,
      Q => blk00000001_sig00000106
    );
  blk00000001_blk00000025_blk00000029 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff3,
      Q => blk00000001_sig00000105
    );
  blk00000001_blk00000025_blk00000028 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff4,
      Q => blk00000001_sig00000104
    );
  blk00000001_blk00000025_blk00000027 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff5,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig0000010e
    );
  blk00000001_blk00000025_blk00000026 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000025_sig00000ff6,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig00000103
    );
  blk00000001_blk000000b1_blk0000010d : INV
    port map (
      I => blk00000001_blk000000b1_sig0000104e,
      O => blk00000001_blk000000b1_sig00001076
    );
  blk00000001_blk000000b1_blk0000010c : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig0000104e,
      I1 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig00001084
    );
  blk00000001_blk000000b1_blk0000010b : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig0000104f,
      I1 => blk00000001_blk000000b1_sig0000104e,
      I2 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig00001082
    );
  blk00000001_blk000000b1_blk0000010a : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig00001050,
      I1 => blk00000001_blk000000b1_sig0000104e,
      I2 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig00001080
    );
  blk00000001_blk000000b1_blk00000109 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig00001051,
      I1 => blk00000001_blk000000b1_sig0000104e,
      I2 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig0000107e
    );
  blk00000001_blk000000b1_blk00000108 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig00001052,
      I1 => blk00000001_blk000000b1_sig0000104e,
      I2 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig0000107c
    );
  blk00000001_blk000000b1_blk00000107 : LUT6
    generic map(
      INIT => X"AAAA2BAAAAAA0AAA"
    )
    port map (
      I0 => blk00000001_sig00000182,
      I1 => blk00000001_blk000000b1_sig0000104e,
      I2 => blk00000001_sig00000181,
      I3 => blk00000001_blk000000b1_sig0000104f,
      I4 => blk00000001_blk000000b1_sig00001086,
      I5 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig00001075
    );
  blk00000001_blk000000b1_blk00000106 : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig00001051,
      I1 => blk00000001_blk000000b1_sig00001050,
      I2 => blk00000001_blk000000b1_sig00001052,
      O => blk00000001_blk000000b1_sig00001086
    );
  blk00000001_blk000000b1_blk00000105 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => blk00000001_blk000000b1_sig0000104e,
      I1 => blk00000001_sig000000f8,
      I2 => blk00000001_sig00000139,
      O => blk00000001_blk000000b1_sig00001085
    );
  blk00000001_blk000000b1_blk00000104 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001085,
      Q => blk00000001_sig0000015c
    );
  blk00000001_blk000000b1_blk00000103 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig000001a3,
      Q => blk00000001_blk000000b1_sig00001054,
      Q15 => NLW_blk00000001_blk000000b1_blk00000103_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk00000102 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig000001a2,
      Q => blk00000001_blk000000b1_sig00001055,
      Q15 => NLW_blk00000001_blk000000b1_blk00000102_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk00000101 : XORCY
    port map (
      CI => blk00000001_blk000000b1_sig00001083,
      LI => blk00000001_blk000000b1_sig00001084,
      O => blk00000001_blk000000b1_sig0000107b
    );
  blk00000001_blk000000b1_blk00000100 : XORCY
    port map (
      CI => blk00000001_blk000000b1_sig00001081,
      LI => blk00000001_blk000000b1_sig00001082,
      O => blk00000001_blk000000b1_sig0000107a
    );
  blk00000001_blk000000b1_blk000000ff : MUXCY
    port map (
      CI => blk00000001_blk000000b1_sig00001081,
      DI => blk00000001_blk000000b1_sig0000104f,
      S => blk00000001_blk000000b1_sig00001082,
      O => blk00000001_blk000000b1_sig00001083
    );
  blk00000001_blk000000b1_blk000000fe : XORCY
    port map (
      CI => blk00000001_blk000000b1_sig0000107f,
      LI => blk00000001_blk000000b1_sig00001080,
      O => blk00000001_blk000000b1_sig00001079
    );
  blk00000001_blk000000b1_blk000000fd : MUXCY
    port map (
      CI => blk00000001_blk000000b1_sig0000107f,
      DI => blk00000001_blk000000b1_sig00001050,
      S => blk00000001_blk000000b1_sig00001080,
      O => blk00000001_blk000000b1_sig00001081
    );
  blk00000001_blk000000b1_blk000000fc : XORCY
    port map (
      CI => blk00000001_blk000000b1_sig0000107d,
      LI => blk00000001_blk000000b1_sig0000107e,
      O => blk00000001_blk000000b1_sig00001078
    );
  blk00000001_blk000000b1_blk000000fb : MUXCY
    port map (
      CI => blk00000001_blk000000b1_sig0000107d,
      DI => blk00000001_blk000000b1_sig00001051,
      S => blk00000001_blk000000b1_sig0000107e,
      O => blk00000001_blk000000b1_sig0000107f
    );
  blk00000001_blk000000b1_blk000000fa : XORCY
    port map (
      CI => blk00000001_sig00000181,
      LI => blk00000001_blk000000b1_sig0000107c,
      O => blk00000001_blk000000b1_sig00001077
    );
  blk00000001_blk000000b1_blk000000f9 : MUXCY
    port map (
      CI => blk00000001_sig00000181,
      DI => blk00000001_blk000000b1_sig00001052,
      S => blk00000001_blk000000b1_sig0000107c,
      O => blk00000001_blk000000b1_sig0000107d
    );
  blk00000001_blk000000b1_blk000000f8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig000001a0,
      Q => blk00000001_blk000000b1_sig00001057,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f8_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019f,
      Q => blk00000001_blk000000b1_sig00001058,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f7_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig000001a1,
      Q => blk00000001_blk000000b1_sig00001056,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f6_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019d,
      Q => blk00000001_blk000000b1_sig0000105a,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f5_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019c,
      Q => blk00000001_blk000000b1_sig0000105b,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f4_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019e,
      Q => blk00000001_blk000000b1_sig00001059,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f3_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019b,
      Q => blk00000001_blk000000b1_sig0000105c,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f2_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000019a,
      Q => blk00000001_blk000000b1_sig0000105d,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f1_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000f0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000199,
      Q => blk00000001_blk000000b1_sig0000105e,
      Q15 => NLW_blk00000001_blk000000b1_blk000000f0_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000ef : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000198,
      Q => blk00000001_blk000000b1_sig0000105f,
      Q15 => NLW_blk00000001_blk000000b1_blk000000ef_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000ee : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000196,
      Q => blk00000001_blk000000b1_sig00001061,
      Q15 => NLW_blk00000001_blk000000b1_blk000000ee_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000ed : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000195,
      Q => blk00000001_blk000000b1_sig00001062,
      Q15 => NLW_blk00000001_blk000000b1_blk000000ed_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000ec : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000197,
      Q => blk00000001_blk000000b1_sig00001060,
      Q15 => NLW_blk00000001_blk000000b1_blk000000ec_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000eb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000193,
      Q => blk00000001_blk000000b1_sig00001064,
      Q15 => NLW_blk00000001_blk000000b1_blk000000eb_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000ea : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000192,
      Q => blk00000001_blk000000b1_sig00001065,
      Q15 => NLW_blk00000001_blk000000b1_blk000000ea_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000194,
      Q => blk00000001_blk000000b1_sig00001063,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e9_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000190,
      Q => blk00000001_blk000000b1_sig00001067,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e8_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018f,
      Q => blk00000001_blk000000b1_sig00001068,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e7_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000191,
      Q => blk00000001_blk000000b1_sig00001066,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e6_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018e,
      Q => blk00000001_blk000000b1_sig00001069,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e5_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018d,
      Q => blk00000001_blk000000b1_sig0000106a,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e4_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018c,
      Q => blk00000001_blk000000b1_sig0000106b,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e3_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018b,
      Q => blk00000001_blk000000b1_sig0000106c,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e2_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000189,
      Q => blk00000001_blk000000b1_sig0000106e,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e1_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000e0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000188,
      Q => blk00000001_blk000000b1_sig0000106f,
      Q15 => NLW_blk00000001_blk000000b1_blk000000e0_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000df : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig0000018a,
      Q => blk00000001_blk000000b1_sig0000106d,
      Q15 => NLW_blk00000001_blk000000b1_blk000000df_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000de : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000186,
      Q => blk00000001_blk000000b1_sig00001071,
      Q15 => NLW_blk00000001_blk000000b1_blk000000de_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000dd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000185,
      Q => blk00000001_blk000000b1_sig00001072,
      Q15 => NLW_blk00000001_blk000000b1_blk000000dd_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000dc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000187,
      Q => blk00000001_blk000000b1_sig00001070,
      Q15 => NLW_blk00000001_blk000000b1_blk000000dc_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000db : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000183,
      Q => blk00000001_blk000000b1_sig00001074,
      Q15 => NLW_blk00000001_blk000000b1_blk000000db_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000da : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000b1_sig00001052,
      A1 => blk00000001_blk000000b1_sig00001051,
      A2 => blk00000001_blk000000b1_sig00001050,
      A3 => blk00000001_blk000000b1_sig0000104f,
      CE => blk00000001_sig00000181,
      CLK => aclk,
      D => blk00000001_sig00000184,
      Q => blk00000001_blk000000b1_sig00001073,
      Q15 => NLW_blk00000001_blk000000b1_blk000000da_Q15_UNCONNECTED
    );
  blk00000001_blk000000b1_blk000000d9 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000107b,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk000000b1_sig0000104e
    );
  blk00000001_blk000000b1_blk000000d8 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000107a,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk000000b1_sig0000104f
    );
  blk00000001_blk000000b1_blk000000d7 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001079,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk000000b1_sig00001050
    );
  blk00000001_blk000000b1_blk000000d6 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001078,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk000000b1_sig00001051
    );
  blk00000001_blk000000b1_blk000000d5 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001077,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk000000b1_sig00001052
    );
  blk00000001_blk000000b1_blk000000d4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001054,
      Q => blk00000001_sig0000017e
    );
  blk00000001_blk000000b1_blk000000d3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001055,
      Q => blk00000001_sig0000017d
    );
  blk00000001_blk000000b1_blk000000d2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001056,
      Q => blk00000001_sig0000017c
    );
  blk00000001_blk000000b1_blk000000d1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001057,
      Q => blk00000001_sig0000017b
    );
  blk00000001_blk000000b1_blk000000d0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001058,
      Q => blk00000001_sig0000017a
    );
  blk00000001_blk000000b1_blk000000cf : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001059,
      Q => blk00000001_sig00000179
    );
  blk00000001_blk000000b1_blk000000ce : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105a,
      Q => blk00000001_sig00000178
    );
  blk00000001_blk000000b1_blk000000cd : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105b,
      Q => blk00000001_sig00000177
    );
  blk00000001_blk000000b1_blk000000cc : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105c,
      Q => blk00000001_sig00000176
    );
  blk00000001_blk000000b1_blk000000cb : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105d,
      Q => blk00000001_sig00000175
    );
  blk00000001_blk000000b1_blk000000ca : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105e,
      Q => blk00000001_sig00000174
    );
  blk00000001_blk000000b1_blk000000c9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000105f,
      Q => blk00000001_sig00000173
    );
  blk00000001_blk000000b1_blk000000c8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001060,
      Q => blk00000001_sig00000172
    );
  blk00000001_blk000000b1_blk000000c7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001061,
      Q => blk00000001_sig00000171
    );
  blk00000001_blk000000b1_blk000000c6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001062,
      Q => blk00000001_sig00000170
    );
  blk00000001_blk000000b1_blk000000c5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001063,
      Q => blk00000001_sig0000016f
    );
  blk00000001_blk000000b1_blk000000c4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001064,
      Q => blk00000001_sig0000016e
    );
  blk00000001_blk000000b1_blk000000c3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001065,
      Q => blk00000001_sig0000016d
    );
  blk00000001_blk000000b1_blk000000c2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001066,
      Q => blk00000001_sig0000016c
    );
  blk00000001_blk000000b1_blk000000c1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001067,
      Q => blk00000001_sig0000016b
    );
  blk00000001_blk000000b1_blk000000c0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001068,
      Q => blk00000001_sig0000016a
    );
  blk00000001_blk000000b1_blk000000bf : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001069,
      Q => blk00000001_sig00000169
    );
  blk00000001_blk000000b1_blk000000be : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106a,
      Q => blk00000001_sig00000168
    );
  blk00000001_blk000000b1_blk000000bd : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106b,
      Q => blk00000001_sig00000167
    );
  blk00000001_blk000000b1_blk000000bc : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106c,
      Q => blk00000001_sig00000166
    );
  blk00000001_blk000000b1_blk000000bb : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106d,
      Q => blk00000001_sig00000165
    );
  blk00000001_blk000000b1_blk000000ba : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106e,
      Q => blk00000001_sig00000164
    );
  blk00000001_blk000000b1_blk000000b9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig0000106f,
      Q => blk00000001_sig00000163
    );
  blk00000001_blk000000b1_blk000000b8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001070,
      Q => blk00000001_sig00000162
    );
  blk00000001_blk000000b1_blk000000b7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001071,
      Q => blk00000001_sig00000161
    );
  blk00000001_blk000000b1_blk000000b6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001072,
      Q => blk00000001_sig00000160
    );
  blk00000001_blk000000b1_blk000000b5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001073,
      Q => blk00000001_sig0000015f
    );
  blk00000001_blk000000b1_blk000000b4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001074,
      Q => blk00000001_sig0000015e
    );
  blk00000001_blk000000b1_blk000000b3 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001075,
      S => blk00000001_sig000000f8,
      Q => blk00000001_sig00000182
    );
  blk00000001_blk000000b1_blk000000b2 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000b1_sig00001076,
      R => blk00000001_sig000000f8,
      Q => blk00000001_sig0000015d
    );
  blk00000001_blk0000010e_blk0000012a : LUT5
    generic map(
      INIT => X"04445544"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      I3 => aclken,
      I4 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig00001096
    );
  blk00000001_blk0000010e_blk00000129 : LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      I3 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig00001097
    );
  blk00000001_blk0000010e_blk00000128 : LUT6
    generic map(
      INIT => X"4044404440444054"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => blk00000001_sig00000100,
      I2 => blk00000001_sig000000d8,
      I3 => blk00000001_blk0000010e_sig000010a6,
      I4 => blk00000001_blk0000010e_sig00001092,
      I5 => blk00000001_blk0000010e_sig000010a8,
      O => blk00000001_blk0000010e_sig000010a7
    );
  blk00000001_blk0000010e_blk00000127 : LUT3
    generic map(
      INIT => X"7F"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig00001091,
      I1 => blk00000001_blk0000010e_sig00001090,
      I2 => blk00000001_blk0000010e_sig0000108f,
      O => blk00000001_blk0000010e_sig000010a8
    );
  blk00000001_blk0000010e_blk00000126 : LUT4
    generic map(
      INIT => X"4044"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig0000108e,
      I1 => aclken,
      I2 => m_axis_status_tready,
      I3 => NlwRenamedSig_OI_m_axis_status_tvalid,
      O => blk00000001_blk0000010e_sig000010a6
    );
  blk00000001_blk0000010e_blk00000125 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig0000108f,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig00001099
    );
  blk00000001_blk0000010e_blk00000124 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig00001090,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig0000109b
    );
  blk00000001_blk0000010e_blk00000123 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig00001091,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig0000109d
    );
  blk00000001_blk0000010e_blk00000122 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000010e_sig00001092,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk0000010e_sig0000108e,
      O => blk00000001_blk0000010e_sig0000109f
    );
  blk00000001_blk0000010e_blk00000121 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a7,
      Q => blk00000001_sig00000100
    );
  blk00000001_blk0000010e_blk00000120 : LUT3
    generic map(
      INIT => X"A2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      O => blk00000001_blk0000010e_sig00001095
    );
  blk00000001_blk0000010e_blk0000011f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000010e_sig00001095,
      D => blk00000001_blk0000010e_sig000010a5,
      Q => m_axis_status_tdata(0)
    );
  blk00000001_blk0000010e_blk0000011e : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a4,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000010e_sig00001092
    );
  blk00000001_blk0000010e_blk0000011d : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a3,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000010e_sig00001091
    );
  blk00000001_blk0000010e_blk0000011c : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a2,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000010e_sig00001090
    );
  blk00000001_blk0000010e_blk0000011b : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a1,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000010e_sig0000108f
    );
  blk00000001_blk0000010e_blk0000011a : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig000010a0,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000010e_sig0000108e
    );
  blk00000001_blk0000010e_blk00000119 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000010e_sig00001092,
      A1 => blk00000001_blk0000010e_sig00001091,
      A2 => blk00000001_blk0000010e_sig00001090,
      A3 => blk00000001_blk0000010e_sig0000108f,
      CE => blk00000001_sig000000d8,
      CLK => aclk,
      D => blk00000001_sig000000f6,
      Q => blk00000001_blk0000010e_sig000010a5,
      Q15 => NLW_blk00000001_blk0000010e_blk00000119_Q15_UNCONNECTED
    );
  blk00000001_blk0000010e_blk00000118 : MUXCY
    port map (
      CI => blk00000001_sig000000d8,
      DI => blk00000001_blk0000010e_sig00001092,
      S => blk00000001_blk0000010e_sig0000109f,
      O => blk00000001_blk0000010e_sig0000109e
    );
  blk00000001_blk0000010e_blk00000117 : XORCY
    port map (
      CI => blk00000001_sig000000d8,
      LI => blk00000001_blk0000010e_sig0000109f,
      O => blk00000001_blk0000010e_sig000010a4
    );
  blk00000001_blk0000010e_blk00000116 : MUXCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109e,
      DI => blk00000001_blk0000010e_sig00001091,
      S => blk00000001_blk0000010e_sig0000109d,
      O => blk00000001_blk0000010e_sig0000109c
    );
  blk00000001_blk0000010e_blk00000115 : XORCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109e,
      LI => blk00000001_blk0000010e_sig0000109d,
      O => blk00000001_blk0000010e_sig000010a3
    );
  blk00000001_blk0000010e_blk00000114 : MUXCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109c,
      DI => blk00000001_blk0000010e_sig00001090,
      S => blk00000001_blk0000010e_sig0000109b,
      O => blk00000001_blk0000010e_sig0000109a
    );
  blk00000001_blk0000010e_blk00000113 : XORCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109c,
      LI => blk00000001_blk0000010e_sig0000109b,
      O => blk00000001_blk0000010e_sig000010a2
    );
  blk00000001_blk0000010e_blk00000112 : MUXCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109a,
      DI => blk00000001_blk0000010e_sig0000108f,
      S => blk00000001_blk0000010e_sig00001099,
      O => blk00000001_blk0000010e_sig00001098
    );
  blk00000001_blk0000010e_blk00000111 : XORCY
    port map (
      CI => blk00000001_blk0000010e_sig0000109a,
      LI => blk00000001_blk0000010e_sig00001099,
      O => blk00000001_blk0000010e_sig000010a1
    );
  blk00000001_blk0000010e_blk00000110 : XORCY
    port map (
      CI => blk00000001_blk0000010e_sig00001098,
      LI => blk00000001_blk0000010e_sig00001097,
      O => blk00000001_blk0000010e_sig000010a0
    );
  blk00000001_blk0000010e_blk0000010f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000010e_sig00001096,
      Q => NlwRenamedSig_OI_m_axis_status_tvalid
    );
  blk00000001_blk0000012b_blk00000198 : LUT5
    generic map(
      INIT => X"04445544"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      I3 => aclken,
      I4 => blk00000001_blk0000012b_sig000010fe,
      O => blk00000001_blk0000012b_sig00001107
    );
  blk00000001_blk0000012b_blk00000197 : LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      I3 => blk00000001_blk0000012b_sig000010fe,
      O => blk00000001_blk0000012b_sig00001108
    );
  blk00000001_blk0000012b_blk00000196 : LUT6
    generic map(
      INIT => X"0A0A0A0B000A000A"
    )
    port map (
      I0 => blk00000001_sig000000ff,
      I1 => blk00000001_blk0000012b_sig00001102,
      I2 => blk00000001_sig000000f8,
      I3 => blk00000001_blk0000012b_sig0000113f,
      I4 => blk00000001_blk0000012b_sig00001142,
      I5 => blk00000001_sig000000da,
      O => blk00000001_blk0000012b_sig00001140
    );
  blk00000001_blk0000012b_blk00000195 : LUT3
    generic map(
      INIT => X"7F"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig00001101,
      I1 => blk00000001_blk0000012b_sig00001100,
      I2 => blk00000001_blk0000012b_sig000010ff,
      O => blk00000001_blk0000012b_sig00001142
    );
  blk00000001_blk0000012b_blk00000194 : LUT4
    generic map(
      INIT => X"4044"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig000010fe,
      I1 => aclken,
      I2 => m_axis_data_tready,
      I3 => NlwRenamedSig_OI_m_axis_data_tvalid,
      O => blk00000001_blk0000012b_sig0000113f
    );
  blk00000001_blk0000012b_blk00000193 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig000010ff,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk0000012b_sig000010fe,
      O => blk00000001_blk0000012b_sig0000110a
    );
  blk00000001_blk0000012b_blk00000192 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig00001100,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk0000012b_sig000010fe,
      O => blk00000001_blk0000012b_sig0000110c
    );
  blk00000001_blk0000012b_blk00000191 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig00001101,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk0000012b_sig000010fe,
      O => blk00000001_blk0000012b_sig0000110e
    );
  blk00000001_blk0000012b_blk00000190 : LUT5
    generic map(
      INIT => X"F7F3080C"
    )
    port map (
      I0 => m_axis_data_tready,
      I1 => aclken,
      I2 => blk00000001_blk0000012b_sig000010fe,
      I3 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I4 => blk00000001_blk0000012b_sig00001102,
      O => blk00000001_blk0000012b_sig00001110
    );
  blk00000001_blk0000012b_blk0000018f : LUT6
    generic map(
      INIT => X"0E0F0A0A080A0A0A"
    )
    port map (
      I0 => blk00000001_sig000000fe,
      I1 => blk00000001_blk0000012b_sig000010fe,
      I2 => blk00000001_sig000000f8,
      I3 => blk00000001_blk0000012b_sig00001106,
      I4 => blk00000001_blk0000012b_sig00001116,
      I5 => blk00000001_sig000000da,
      O => blk00000001_blk0000012b_sig00001141
    );
  blk00000001_blk0000012b_blk0000018e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001141,
      Q => blk00000001_sig000000fe
    );
  blk00000001_blk0000012b_blk0000018d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001140,
      Q => blk00000001_sig000000ff
    );
  blk00000001_blk0000012b_blk0000018c : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => blk00000001_blk0000012b_sig000010ff,
      I1 => blk00000001_blk0000012b_sig00001100,
      I2 => blk00000001_blk0000012b_sig00001101,
      I3 => blk00000001_blk0000012b_sig00001102,
      O => blk00000001_blk0000012b_sig00001116
    );
  blk00000001_blk0000012b_blk0000018b : LUT3
    generic map(
      INIT => X"A2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      O => blk00000001_blk0000012b_sig00001106
    );
  blk00000001_blk0000012b_blk0000018a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001117,
      Q => m_axis_data_tlast
    );
  blk00000001_blk0000012b_blk00000189 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001118,
      Q => m_axis_data_tdata(0)
    );
  blk00000001_blk0000012b_blk00000188 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001119,
      Q => m_axis_data_tdata(1)
    );
  blk00000001_blk0000012b_blk00000187 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111a,
      Q => m_axis_data_tdata(2)
    );
  blk00000001_blk0000012b_blk00000186 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111b,
      Q => m_axis_data_tdata(3)
    );
  blk00000001_blk0000012b_blk00000185 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111c,
      Q => m_axis_data_tdata(4)
    );
  blk00000001_blk0000012b_blk00000184 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111d,
      Q => m_axis_data_tdata(5)
    );
  blk00000001_blk0000012b_blk00000183 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111e,
      Q => m_axis_data_tdata(6)
    );
  blk00000001_blk0000012b_blk00000182 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000111f,
      Q => m_axis_data_tdata(7)
    );
  blk00000001_blk0000012b_blk00000181 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001120,
      Q => m_axis_data_tdata(8)
    );
  blk00000001_blk0000012b_blk00000180 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001121,
      Q => m_axis_data_tdata(9)
    );
  blk00000001_blk0000012b_blk0000017f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001122,
      Q => m_axis_data_tdata(10)
    );
  blk00000001_blk0000012b_blk0000017e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001123,
      Q => m_axis_data_tdata(11)
    );
  blk00000001_blk0000012b_blk0000017d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001124,
      Q => m_axis_data_tdata(12)
    );
  blk00000001_blk0000012b_blk0000017c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001125,
      Q => m_axis_data_tdata(13)
    );
  blk00000001_blk0000012b_blk0000017b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001126,
      Q => m_axis_data_tdata(14)
    );
  blk00000001_blk0000012b_blk0000017a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001127,
      Q => m_axis_data_tdata(15)
    );
  blk00000001_blk0000012b_blk00000179 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001128,
      Q => m_axis_data_tdata(16)
    );
  blk00000001_blk0000012b_blk00000178 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001129,
      Q => m_axis_data_tdata(17)
    );
  blk00000001_blk0000012b_blk00000177 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112a,
      Q => m_axis_data_tdata(18)
    );
  blk00000001_blk0000012b_blk00000176 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112b,
      Q => m_axis_data_tdata(19)
    );
  blk00000001_blk0000012b_blk00000175 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112c,
      Q => m_axis_data_tdata(20)
    );
  blk00000001_blk0000012b_blk00000174 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112d,
      Q => m_axis_data_tdata(21)
    );
  blk00000001_blk0000012b_blk00000173 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112e,
      Q => m_axis_data_tdata(22)
    );
  blk00000001_blk0000012b_blk00000172 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000112f,
      Q => m_axis_data_tdata(23)
    );
  blk00000001_blk0000012b_blk00000171 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001130,
      Q => m_axis_data_tdata(24)
    );
  blk00000001_blk0000012b_blk00000170 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001131,
      Q => m_axis_data_tdata(25)
    );
  blk00000001_blk0000012b_blk0000016f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001132,
      Q => m_axis_data_tdata(26)
    );
  blk00000001_blk0000012b_blk0000016e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001133,
      Q => m_axis_data_tdata(27)
    );
  blk00000001_blk0000012b_blk0000016d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001134,
      Q => m_axis_data_tdata(28)
    );
  blk00000001_blk0000012b_blk0000016c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001135,
      Q => m_axis_data_tdata(29)
    );
  blk00000001_blk0000012b_blk0000016b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001136,
      Q => m_axis_data_tdata(30)
    );
  blk00000001_blk0000012b_blk0000016a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001137,
      Q => m_axis_data_tdata(31)
    );
  blk00000001_blk0000012b_blk00000169 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001138,
      Q => m_axis_data_tuser(0)
    );
  blk00000001_blk0000012b_blk00000168 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig00001139,
      Q => m_axis_data_tuser(1)
    );
  blk00000001_blk0000012b_blk00000167 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000113a,
      Q => m_axis_data_tuser(2)
    );
  blk00000001_blk0000012b_blk00000166 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000113b,
      Q => m_axis_data_tuser(3)
    );
  blk00000001_blk0000012b_blk00000165 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000113c,
      Q => m_axis_data_tuser(4)
    );
  blk00000001_blk0000012b_blk00000164 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000113d,
      Q => m_axis_data_tuser(5)
    );
  blk00000001_blk0000012b_blk00000163 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk0000012b_sig00001106,
      D => blk00000001_blk0000012b_sig0000113e,
      Q => NlwRenamedSig_OI_m_axis_data_tuser_8_Q
    );
  blk00000001_blk0000012b_blk00000162 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001115,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000012b_sig00001102
    );
  blk00000001_blk0000012b_blk00000161 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001114,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000012b_sig00001101
    );
  blk00000001_blk0000012b_blk00000160 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001113,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000012b_sig00001100
    );
  blk00000001_blk0000012b_blk0000015f : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001112,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000012b_sig000010ff
    );
  blk00000001_blk0000012b_blk0000015e : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001111,
      S => blk00000001_sig000000f8,
      Q => blk00000001_blk0000012b_sig000010fe
    );
  blk00000001_blk0000012b_blk0000015d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000db,
      Q => blk00000001_blk0000012b_sig00001117,
      Q15 => NLW_blk00000001_blk0000012b_blk0000015d_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000015c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000aa,
      Q => blk00000001_blk0000012b_sig00001118,
      Q15 => NLW_blk00000001_blk0000012b_blk0000015c_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000015b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a9,
      Q => blk00000001_blk0000012b_sig00001119,
      Q15 => NLW_blk00000001_blk0000012b_blk0000015b_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000015a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a6,
      Q => blk00000001_blk0000012b_sig0000111c,
      Q15 => NLW_blk00000001_blk0000012b_blk0000015a_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000159 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a8,
      Q => blk00000001_blk0000012b_sig0000111a,
      Q15 => NLW_blk00000001_blk0000012b_blk00000159_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000158 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a7,
      Q => blk00000001_blk0000012b_sig0000111b,
      Q15 => NLW_blk00000001_blk0000012b_blk00000158_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000157 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a5,
      Q => blk00000001_blk0000012b_sig0000111d,
      Q15 => NLW_blk00000001_blk0000012b_blk00000157_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000156 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a4,
      Q => blk00000001_blk0000012b_sig0000111e,
      Q15 => NLW_blk00000001_blk0000012b_blk00000156_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000155 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a3,
      Q => blk00000001_blk0000012b_sig0000111f,
      Q15 => NLW_blk00000001_blk0000012b_blk00000155_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000154 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a2,
      Q => blk00000001_blk0000012b_sig00001120,
      Q15 => NLW_blk00000001_blk0000012b_blk00000154_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000153 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009f,
      Q => blk00000001_blk0000012b_sig00001123,
      Q15 => NLW_blk00000001_blk0000012b_blk00000153_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000152 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a1,
      Q => blk00000001_blk0000012b_sig00001121,
      Q15 => NLW_blk00000001_blk0000012b_blk00000152_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000151 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000a0,
      Q => blk00000001_blk0000012b_sig00001122,
      Q15 => NLW_blk00000001_blk0000012b_blk00000151_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000150 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009e,
      Q => blk00000001_blk0000012b_sig00001124,
      Q15 => NLW_blk00000001_blk0000012b_blk00000150_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009d,
      Q => blk00000001_blk0000012b_sig00001125,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014f_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009c,
      Q => blk00000001_blk0000012b_sig00001126,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014e_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009b,
      Q => blk00000001_blk0000012b_sig00001127,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014d_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b8,
      Q => blk00000001_blk0000012b_sig0000112a,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014c_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000ba,
      Q => blk00000001_blk0000012b_sig00001128,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014b_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000014a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b9,
      Q => blk00000001_blk0000012b_sig00001129,
      Q15 => NLW_blk00000001_blk0000012b_blk0000014a_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000149 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b7,
      Q => blk00000001_blk0000012b_sig0000112b,
      Q15 => NLW_blk00000001_blk0000012b_blk00000149_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000148 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b6,
      Q => blk00000001_blk0000012b_sig0000112c,
      Q15 => NLW_blk00000001_blk0000012b_blk00000148_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000147 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b5,
      Q => blk00000001_blk0000012b_sig0000112d,
      Q15 => NLW_blk00000001_blk0000012b_blk00000147_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000146 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b4,
      Q => blk00000001_blk0000012b_sig0000112e,
      Q15 => NLW_blk00000001_blk0000012b_blk00000146_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000145 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b1,
      Q => blk00000001_blk0000012b_sig00001131,
      Q15 => NLW_blk00000001_blk0000012b_blk00000145_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000144 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b3,
      Q => blk00000001_blk0000012b_sig0000112f,
      Q15 => NLW_blk00000001_blk0000012b_blk00000144_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000143 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b2,
      Q => blk00000001_blk0000012b_sig00001130,
      Q15 => NLW_blk00000001_blk0000012b_blk00000143_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000142 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000b0,
      Q => blk00000001_blk0000012b_sig00001132,
      Q15 => NLW_blk00000001_blk0000012b_blk00000142_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000141 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000af,
      Q => blk00000001_blk0000012b_sig00001133,
      Q15 => NLW_blk00000001_blk0000012b_blk00000141_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000140 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000ae,
      Q => blk00000001_blk0000012b_sig00001134,
      Q15 => NLW_blk00000001_blk0000012b_blk00000140_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000ad,
      Q => blk00000001_blk0000012b_sig00001135,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013f_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig0000009a,
      Q => blk00000001_blk0000012b_sig00001138,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013e_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000ac,
      Q => blk00000001_blk0000012b_sig00001136,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013d_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000ab,
      Q => blk00000001_blk0000012b_sig00001137,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013c_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig00000099,
      Q => blk00000001_blk0000012b_sig00001139,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013b_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000013a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig00000098,
      Q => blk00000001_blk0000012b_sig0000113a,
      Q15 => NLW_blk00000001_blk0000012b_blk0000013a_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000139 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig00000097,
      Q => blk00000001_blk0000012b_sig0000113b,
      Q15 => NLW_blk00000001_blk0000012b_blk00000139_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000138 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig00000096,
      Q => blk00000001_blk0000012b_sig0000113c,
      Q15 => NLW_blk00000001_blk0000012b_blk00000138_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk00000137 : MUXCY
    port map (
      CI => blk00000001_sig000000da,
      DI => blk00000001_blk0000012b_sig00001102,
      S => blk00000001_blk0000012b_sig00001110,
      O => blk00000001_blk0000012b_sig0000110f
    );
  blk00000001_blk0000012b_blk00000136 : XORCY
    port map (
      CI => blk00000001_sig000000da,
      LI => blk00000001_blk0000012b_sig00001110,
      O => blk00000001_blk0000012b_sig00001115
    );
  blk00000001_blk0000012b_blk00000135 : MUXCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110f,
      DI => blk00000001_blk0000012b_sig00001101,
      S => blk00000001_blk0000012b_sig0000110e,
      O => blk00000001_blk0000012b_sig0000110d
    );
  blk00000001_blk0000012b_blk00000134 : XORCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110f,
      LI => blk00000001_blk0000012b_sig0000110e,
      O => blk00000001_blk0000012b_sig00001114
    );
  blk00000001_blk0000012b_blk00000133 : MUXCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110d,
      DI => blk00000001_blk0000012b_sig00001100,
      S => blk00000001_blk0000012b_sig0000110c,
      O => blk00000001_blk0000012b_sig0000110b
    );
  blk00000001_blk0000012b_blk00000132 : XORCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110d,
      LI => blk00000001_blk0000012b_sig0000110c,
      O => blk00000001_blk0000012b_sig00001113
    );
  blk00000001_blk0000012b_blk00000131 : MUXCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110b,
      DI => blk00000001_blk0000012b_sig000010ff,
      S => blk00000001_blk0000012b_sig0000110a,
      O => blk00000001_blk0000012b_sig00001109
    );
  blk00000001_blk0000012b_blk00000130 : XORCY
    port map (
      CI => blk00000001_blk0000012b_sig0000110b,
      LI => blk00000001_blk0000012b_sig0000110a,
      O => blk00000001_blk0000012b_sig00001112
    );
  blk00000001_blk0000012b_blk0000012f : XORCY
    port map (
      CI => blk00000001_blk0000012b_sig00001109,
      LI => blk00000001_blk0000012b_sig00001108,
      O => blk00000001_blk0000012b_sig00001111
    );
  blk00000001_blk0000012b_blk0000012e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig00000095,
      Q => blk00000001_blk0000012b_sig0000113d,
      Q15 => NLW_blk00000001_blk0000012b_blk0000012e_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000012d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000012b_sig00001102,
      A1 => blk00000001_blk0000012b_sig00001101,
      A2 => blk00000001_blk0000012b_sig00001100,
      A3 => blk00000001_blk0000012b_sig000010ff,
      CE => blk00000001_sig000000da,
      CLK => aclk,
      D => blk00000001_sig000000bf,
      Q => blk00000001_blk0000012b_sig0000113e,
      Q15 => NLW_blk00000001_blk0000012b_blk0000012d_Q15_UNCONNECTED
    );
  blk00000001_blk0000012b_blk0000012c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk0000012b_sig00001107,
      Q => NlwRenamedSig_OI_m_axis_data_tvalid
    );
  blk00000001_blk000007e0_blk000007e1_blk000007e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000007e0_blk000007e1_sig0000114e,
      Q => blk00000001_sig000002e1
    );
  blk00000001_blk000007e0_blk000007e1_blk000007e4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000007e0_blk000007e1_sig0000114d,
      A1 => blk00000001_blk000007e0_blk000007e1_sig0000114c,
      A2 => blk00000001_blk000007e0_blk000007e1_sig0000114c,
      A3 => blk00000001_blk000007e0_blk000007e1_sig0000114c,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001a6,
      Q => blk00000001_blk000007e0_blk000007e1_sig0000114e,
      Q15 => NLW_blk00000001_blk000007e0_blk000007e1_blk000007e4_Q15_UNCONNECTED
    );
  blk00000001_blk000007e0_blk000007e1_blk000007e3 : VCC
    port map (
      P => blk00000001_blk000007e0_blk000007e1_sig0000114d
    );
  blk00000001_blk000007e0_blk000007e1_blk000007e2 : GND
    port map (
      G => blk00000001_blk000007e0_blk000007e1_sig0000114c
    );
  blk00000001_blk000008e6_blk00000908 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000008e,
      RDCLK => aclk,
      WREN => blk00000001_sig0000008e,
      RDEN => blk00000001_sig0000008e,
      WRCLK => aclk,
      SSR => blk00000001_blk000008e6_sig000011bb,
      DIP(3) => blk00000001_blk000008e6_sig000011bb,
      DIP(2) => blk00000001_sig0000027b,
      DIP(1) => blk00000001_sig00000272,
      DIP(0) => blk00000001_sig00000269,
      DOP(3) => NLW_blk00000001_blk000008e6_blk00000908_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk000008e6_sig0000119a,
      DOP(1) => blk00000001_blk000008e6_sig00001199,
      DOP(0) => blk00000001_blk000008e6_sig00001198,
      WE(3) => blk00000001_sig000001d5,
      WE(2) => blk00000001_sig000001d5,
      WE(1) => blk00000001_sig000001d5,
      WE(0) => blk00000001_sig000001d5,
      DO(31) => NLW_blk00000001_blk000008e6_blk00000908_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk000008e6_blk00000908_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk000008e6_blk00000908_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk000008e6_sig00001193,
      DO(27) => blk00000001_blk000008e6_sig00001194,
      DO(26) => blk00000001_blk000008e6_sig00001195,
      DO(25) => blk00000001_blk000008e6_sig00001196,
      DO(24) => blk00000001_blk000008e6_sig00001197,
      DO(23) => blk00000001_blk000008e6_sig0000118b,
      DO(22) => blk00000001_blk000008e6_sig0000118c,
      DO(21) => blk00000001_blk000008e6_sig0000118d,
      DO(20) => blk00000001_blk000008e6_sig0000118e,
      DO(19) => blk00000001_blk000008e6_sig0000118f,
      DO(18) => blk00000001_blk000008e6_sig00001190,
      DO(17) => blk00000001_blk000008e6_sig00001191,
      DO(16) => blk00000001_blk000008e6_sig00001192,
      DO(15) => blk00000001_blk000008e6_sig00001183,
      DO(14) => blk00000001_blk000008e6_sig00001184,
      DO(13) => blk00000001_blk000008e6_sig00001185,
      DO(12) => blk00000001_blk000008e6_sig00001186,
      DO(11) => blk00000001_blk000008e6_sig00001187,
      DO(10) => blk00000001_blk000008e6_sig00001188,
      DO(9) => blk00000001_blk000008e6_sig00001189,
      DO(8) => blk00000001_blk000008e6_sig0000118a,
      DO(7) => blk00000001_blk000008e6_sig0000117b,
      DO(6) => blk00000001_blk000008e6_sig0000117c,
      DO(5) => blk00000001_blk000008e6_sig0000117d,
      DO(4) => blk00000001_blk000008e6_sig0000117e,
      DO(3) => blk00000001_blk000008e6_sig0000117f,
      DO(2) => blk00000001_blk000008e6_sig00001180,
      DO(1) => blk00000001_blk000008e6_sig00001181,
      DO(0) => blk00000001_blk000008e6_sig00001182,
      WRADDR(8) => blk00000001_sig000001c8,
      WRADDR(7) => blk00000001_sig000001c7,
      WRADDR(6) => blk00000001_sig000001c6,
      WRADDR(5) => blk00000001_sig000001c5,
      WRADDR(4) => blk00000001_blk000008e6_sig000011bb,
      WRADDR(3) => blk00000001_blk000008e6_sig000011bb,
      WRADDR(2) => blk00000001_blk000008e6_sig000011bb,
      WRADDR(1) => blk00000001_blk000008e6_sig000011bb,
      WRADDR(0) => blk00000001_blk000008e6_sig000011bb,
      RDADDR(8) => blk00000001_sig000001bb,
      RDADDR(7) => blk00000001_sig000001bf,
      RDADDR(6) => blk00000001_sig000001ba,
      RDADDR(5) => blk00000001_sig000001b9,
      RDADDR(4) => blk00000001_blk000008e6_sig000011bb,
      RDADDR(3) => blk00000001_blk000008e6_sig000011bb,
      RDADDR(2) => blk00000001_blk000008e6_sig000011bb,
      RDADDR(1) => blk00000001_blk000008e6_sig000011bb,
      RDADDR(0) => blk00000001_blk000008e6_sig000011bb,
      DI(31) => blk00000001_blk000008e6_sig000011bb,
      DI(30) => blk00000001_blk000008e6_sig000011bb,
      DI(29) => blk00000001_blk000008e6_sig000011bb,
      DI(28) => blk00000001_sig00000280,
      DI(27) => blk00000001_sig0000027f,
      DI(26) => blk00000001_sig0000027e,
      DI(25) => blk00000001_sig0000027d,
      DI(24) => blk00000001_sig0000027c,
      DI(23) => blk00000001_sig0000027a,
      DI(22) => blk00000001_sig00000279,
      DI(21) => blk00000001_sig00000278,
      DI(20) => blk00000001_sig00000277,
      DI(19) => blk00000001_sig00000276,
      DI(18) => blk00000001_sig00000275,
      DI(17) => blk00000001_sig00000274,
      DI(16) => blk00000001_sig00000273,
      DI(15) => blk00000001_sig00000271,
      DI(14) => blk00000001_sig00000270,
      DI(13) => blk00000001_sig0000026f,
      DI(12) => blk00000001_sig0000026e,
      DI(11) => blk00000001_sig0000026d,
      DI(10) => blk00000001_sig0000026c,
      DI(9) => blk00000001_sig0000026b,
      DI(8) => blk00000001_sig0000026a,
      DI(7) => blk00000001_sig00000268,
      DI(6) => blk00000001_sig00000267,
      DI(5) => blk00000001_sig00000266,
      DI(4) => blk00000001_sig00000265,
      DI(3) => blk00000001_sig00000264,
      DI(2) => blk00000001_sig00000263,
      DI(1) => blk00000001_sig00000262,
      DI(0) => blk00000001_sig00000261
    );
  blk00000001_blk000008e6_blk00000907 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001193,
      Q => blk00000001_sig00000200
    );
  blk00000001_blk000008e6_blk00000906 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001194,
      Q => blk00000001_sig000001ff
    );
  blk00000001_blk000008e6_blk00000905 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001195,
      Q => blk00000001_sig000001fe
    );
  blk00000001_blk000008e6_blk00000904 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001196,
      Q => blk00000001_sig000001fd
    );
  blk00000001_blk000008e6_blk00000903 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001197,
      Q => blk00000001_sig000001fc
    );
  blk00000001_blk000008e6_blk00000902 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000119a,
      Q => blk00000001_sig000001fb
    );
  blk00000001_blk000008e6_blk00000901 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118b,
      Q => blk00000001_sig000001fa
    );
  blk00000001_blk000008e6_blk00000900 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118c,
      Q => blk00000001_sig000001f9
    );
  blk00000001_blk000008e6_blk000008ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118d,
      Q => blk00000001_sig000001f8
    );
  blk00000001_blk000008e6_blk000008fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118e,
      Q => blk00000001_sig000001f7
    );
  blk00000001_blk000008e6_blk000008fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118f,
      Q => blk00000001_sig000001f6
    );
  blk00000001_blk000008e6_blk000008fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001190,
      Q => blk00000001_sig000001f5
    );
  blk00000001_blk000008e6_blk000008fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001191,
      Q => blk00000001_sig000001f4
    );
  blk00000001_blk000008e6_blk000008fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001192,
      Q => blk00000001_sig000001f3
    );
  blk00000001_blk000008e6_blk000008f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001199,
      Q => blk00000001_sig000001f2
    );
  blk00000001_blk000008e6_blk000008f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001183,
      Q => blk00000001_sig000001f1
    );
  blk00000001_blk000008e6_blk000008f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001184,
      Q => blk00000001_sig000001f0
    );
  blk00000001_blk000008e6_blk000008f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001185,
      Q => blk00000001_sig000001ef
    );
  blk00000001_blk000008e6_blk000008f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001186,
      Q => blk00000001_sig000001ee
    );
  blk00000001_blk000008e6_blk000008f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001187,
      Q => blk00000001_sig000001ed
    );
  blk00000001_blk000008e6_blk000008f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001188,
      Q => blk00000001_sig000001ec
    );
  blk00000001_blk000008e6_blk000008f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001189,
      Q => blk00000001_sig000001eb
    );
  blk00000001_blk000008e6_blk000008f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000118a,
      Q => blk00000001_sig000001ea
    );
  blk00000001_blk000008e6_blk000008f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001198,
      Q => blk00000001_sig000001e9
    );
  blk00000001_blk000008e6_blk000008ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000117b,
      Q => blk00000001_sig000001e8
    );
  blk00000001_blk000008e6_blk000008ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000117c,
      Q => blk00000001_sig000001e7
    );
  blk00000001_blk000008e6_blk000008ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000117d,
      Q => blk00000001_sig000001e6
    );
  blk00000001_blk000008e6_blk000008ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000117e,
      Q => blk00000001_sig000001e5
    );
  blk00000001_blk000008e6_blk000008eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig0000117f,
      Q => blk00000001_sig000001e4
    );
  blk00000001_blk000008e6_blk000008ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001180,
      Q => blk00000001_sig000001e3
    );
  blk00000001_blk000008e6_blk000008e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001181,
      Q => blk00000001_sig000001e2
    );
  blk00000001_blk000008e6_blk000008e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk000008e6_sig00001182,
      Q => blk00000001_sig000001e1
    );
  blk00000001_blk000008e6_blk000008e7 : GND
    port map (
      G => blk00000001_blk000008e6_sig000011bb
    );
  blk00000001_blk00000909_blk0000092b : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000008e,
      RDCLK => aclk,
      WREN => blk00000001_sig0000008e,
      RDEN => blk00000001_sig0000008e,
      WRCLK => aclk,
      SSR => blk00000001_blk00000909_sig00001228,
      DIP(3) => blk00000001_blk00000909_sig00001228,
      DIP(2) => blk00000001_sig0000029b,
      DIP(1) => blk00000001_sig00000292,
      DIP(0) => blk00000001_sig00000289,
      DOP(3) => NLW_blk00000001_blk00000909_blk0000092b_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk00000909_sig00001207,
      DOP(1) => blk00000001_blk00000909_sig00001206,
      DOP(0) => blk00000001_blk00000909_sig00001205,
      WE(3) => blk00000001_sig000001d6,
      WE(2) => blk00000001_sig000001d6,
      WE(1) => blk00000001_sig000001d6,
      WE(0) => blk00000001_sig000001d6,
      DO(31) => NLW_blk00000001_blk00000909_blk0000092b_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk00000909_blk0000092b_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk00000909_blk0000092b_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk00000909_sig00001200,
      DO(27) => blk00000001_blk00000909_sig00001201,
      DO(26) => blk00000001_blk00000909_sig00001202,
      DO(25) => blk00000001_blk00000909_sig00001203,
      DO(24) => blk00000001_blk00000909_sig00001204,
      DO(23) => blk00000001_blk00000909_sig000011f8,
      DO(22) => blk00000001_blk00000909_sig000011f9,
      DO(21) => blk00000001_blk00000909_sig000011fa,
      DO(20) => blk00000001_blk00000909_sig000011fb,
      DO(19) => blk00000001_blk00000909_sig000011fc,
      DO(18) => blk00000001_blk00000909_sig000011fd,
      DO(17) => blk00000001_blk00000909_sig000011fe,
      DO(16) => blk00000001_blk00000909_sig000011ff,
      DO(15) => blk00000001_blk00000909_sig000011f0,
      DO(14) => blk00000001_blk00000909_sig000011f1,
      DO(13) => blk00000001_blk00000909_sig000011f2,
      DO(12) => blk00000001_blk00000909_sig000011f3,
      DO(11) => blk00000001_blk00000909_sig000011f4,
      DO(10) => blk00000001_blk00000909_sig000011f5,
      DO(9) => blk00000001_blk00000909_sig000011f6,
      DO(8) => blk00000001_blk00000909_sig000011f7,
      DO(7) => blk00000001_blk00000909_sig000011e8,
      DO(6) => blk00000001_blk00000909_sig000011e9,
      DO(5) => blk00000001_blk00000909_sig000011ea,
      DO(4) => blk00000001_blk00000909_sig000011eb,
      DO(3) => blk00000001_blk00000909_sig000011ec,
      DO(2) => blk00000001_blk00000909_sig000011ed,
      DO(1) => blk00000001_blk00000909_sig000011ee,
      DO(0) => blk00000001_blk00000909_sig000011ef,
      WRADDR(8) => blk00000001_sig000001cc,
      WRADDR(7) => blk00000001_sig000001cb,
      WRADDR(6) => blk00000001_sig000001ca,
      WRADDR(5) => blk00000001_sig000001c9,
      WRADDR(4) => blk00000001_blk00000909_sig00001228,
      WRADDR(3) => blk00000001_blk00000909_sig00001228,
      WRADDR(2) => blk00000001_blk00000909_sig00001228,
      WRADDR(1) => blk00000001_blk00000909_sig00001228,
      WRADDR(0) => blk00000001_blk00000909_sig00001228,
      RDADDR(8) => blk00000001_sig000001bd,
      RDADDR(7) => blk00000001_sig000001c3,
      RDADDR(6) => blk00000001_sig000001bc,
      RDADDR(5) => blk00000001_sig000001c1,
      RDADDR(4) => blk00000001_blk00000909_sig00001228,
      RDADDR(3) => blk00000001_blk00000909_sig00001228,
      RDADDR(2) => blk00000001_blk00000909_sig00001228,
      RDADDR(1) => blk00000001_blk00000909_sig00001228,
      RDADDR(0) => blk00000001_blk00000909_sig00001228,
      DI(31) => blk00000001_blk00000909_sig00001228,
      DI(30) => blk00000001_blk00000909_sig00001228,
      DI(29) => blk00000001_blk00000909_sig00001228,
      DI(28) => blk00000001_sig000002a0,
      DI(27) => blk00000001_sig0000029f,
      DI(26) => blk00000001_sig0000029e,
      DI(25) => blk00000001_sig0000029d,
      DI(24) => blk00000001_sig0000029c,
      DI(23) => blk00000001_sig0000029a,
      DI(22) => blk00000001_sig00000299,
      DI(21) => blk00000001_sig00000298,
      DI(20) => blk00000001_sig00000297,
      DI(19) => blk00000001_sig00000296,
      DI(18) => blk00000001_sig00000295,
      DI(17) => blk00000001_sig00000294,
      DI(16) => blk00000001_sig00000293,
      DI(15) => blk00000001_sig00000291,
      DI(14) => blk00000001_sig00000290,
      DI(13) => blk00000001_sig0000028f,
      DI(12) => blk00000001_sig0000028e,
      DI(11) => blk00000001_sig0000028d,
      DI(10) => blk00000001_sig0000028c,
      DI(9) => blk00000001_sig0000028b,
      DI(8) => blk00000001_sig0000028a,
      DI(7) => blk00000001_sig00000288,
      DI(6) => blk00000001_sig00000287,
      DI(5) => blk00000001_sig00000286,
      DI(4) => blk00000001_sig00000285,
      DI(3) => blk00000001_sig00000284,
      DI(2) => blk00000001_sig00000283,
      DI(1) => blk00000001_sig00000282,
      DI(0) => blk00000001_sig00000281
    );
  blk00000001_blk00000909_blk0000092a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001200,
      Q => blk00000001_sig00000220
    );
  blk00000001_blk00000909_blk00000929 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001201,
      Q => blk00000001_sig0000021f
    );
  blk00000001_blk00000909_blk00000928 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001202,
      Q => blk00000001_sig0000021e
    );
  blk00000001_blk00000909_blk00000927 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001203,
      Q => blk00000001_sig0000021d
    );
  blk00000001_blk00000909_blk00000926 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001204,
      Q => blk00000001_sig0000021c
    );
  blk00000001_blk00000909_blk00000925 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001207,
      Q => blk00000001_sig0000021b
    );
  blk00000001_blk00000909_blk00000924 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f8,
      Q => blk00000001_sig0000021a
    );
  blk00000001_blk00000909_blk00000923 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f9,
      Q => blk00000001_sig00000219
    );
  blk00000001_blk00000909_blk00000922 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011fa,
      Q => blk00000001_sig00000218
    );
  blk00000001_blk00000909_blk00000921 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011fb,
      Q => blk00000001_sig00000217
    );
  blk00000001_blk00000909_blk00000920 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011fc,
      Q => blk00000001_sig00000216
    );
  blk00000001_blk00000909_blk0000091f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011fd,
      Q => blk00000001_sig00000215
    );
  blk00000001_blk00000909_blk0000091e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011fe,
      Q => blk00000001_sig00000214
    );
  blk00000001_blk00000909_blk0000091d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ff,
      Q => blk00000001_sig00000213
    );
  blk00000001_blk00000909_blk0000091c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001206,
      Q => blk00000001_sig00000212
    );
  blk00000001_blk00000909_blk0000091b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f0,
      Q => blk00000001_sig00000211
    );
  blk00000001_blk00000909_blk0000091a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f1,
      Q => blk00000001_sig00000210
    );
  blk00000001_blk00000909_blk00000919 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f2,
      Q => blk00000001_sig0000020f
    );
  blk00000001_blk00000909_blk00000918 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f3,
      Q => blk00000001_sig0000020e
    );
  blk00000001_blk00000909_blk00000917 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f4,
      Q => blk00000001_sig0000020d
    );
  blk00000001_blk00000909_blk00000916 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f5,
      Q => blk00000001_sig0000020c
    );
  blk00000001_blk00000909_blk00000915 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f6,
      Q => blk00000001_sig0000020b
    );
  blk00000001_blk00000909_blk00000914 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011f7,
      Q => blk00000001_sig0000020a
    );
  blk00000001_blk00000909_blk00000913 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig00001205,
      Q => blk00000001_sig00000209
    );
  blk00000001_blk00000909_blk00000912 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011e8,
      Q => blk00000001_sig00000208
    );
  blk00000001_blk00000909_blk00000911 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011e9,
      Q => blk00000001_sig00000207
    );
  blk00000001_blk00000909_blk00000910 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ea,
      Q => blk00000001_sig00000206
    );
  blk00000001_blk00000909_blk0000090f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011eb,
      Q => blk00000001_sig00000205
    );
  blk00000001_blk00000909_blk0000090e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ec,
      Q => blk00000001_sig00000204
    );
  blk00000001_blk00000909_blk0000090d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ed,
      Q => blk00000001_sig00000203
    );
  blk00000001_blk00000909_blk0000090c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ee,
      Q => blk00000001_sig00000202
    );
  blk00000001_blk00000909_blk0000090b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000909_sig000011ef,
      Q => blk00000001_sig00000201
    );
  blk00000001_blk00000909_blk0000090a : GND
    port map (
      G => blk00000001_blk00000909_sig00001228
    );
  blk00000001_blk0000092c_blk0000094e : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000008e,
      RDCLK => aclk,
      WREN => blk00000001_sig0000008e,
      RDEN => blk00000001_sig0000008e,
      WRCLK => aclk,
      SSR => blk00000001_blk0000092c_sig00001295,
      DIP(3) => blk00000001_blk0000092c_sig00001295,
      DIP(2) => blk00000001_sig000002bb,
      DIP(1) => blk00000001_sig000002b2,
      DIP(0) => blk00000001_sig000002a9,
      DOP(3) => NLW_blk00000001_blk0000092c_blk0000094e_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk0000092c_sig00001274,
      DOP(1) => blk00000001_blk0000092c_sig00001273,
      DOP(0) => blk00000001_blk0000092c_sig00001272,
      WE(3) => blk00000001_sig000001d7,
      WE(2) => blk00000001_sig000001d7,
      WE(1) => blk00000001_sig000001d7,
      WE(0) => blk00000001_sig000001d7,
      DO(31) => NLW_blk00000001_blk0000092c_blk0000094e_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk0000092c_blk0000094e_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk0000092c_blk0000094e_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk0000092c_sig0000126d,
      DO(27) => blk00000001_blk0000092c_sig0000126e,
      DO(26) => blk00000001_blk0000092c_sig0000126f,
      DO(25) => blk00000001_blk0000092c_sig00001270,
      DO(24) => blk00000001_blk0000092c_sig00001271,
      DO(23) => blk00000001_blk0000092c_sig00001265,
      DO(22) => blk00000001_blk0000092c_sig00001266,
      DO(21) => blk00000001_blk0000092c_sig00001267,
      DO(20) => blk00000001_blk0000092c_sig00001268,
      DO(19) => blk00000001_blk0000092c_sig00001269,
      DO(18) => blk00000001_blk0000092c_sig0000126a,
      DO(17) => blk00000001_blk0000092c_sig0000126b,
      DO(16) => blk00000001_blk0000092c_sig0000126c,
      DO(15) => blk00000001_blk0000092c_sig0000125d,
      DO(14) => blk00000001_blk0000092c_sig0000125e,
      DO(13) => blk00000001_blk0000092c_sig0000125f,
      DO(12) => blk00000001_blk0000092c_sig00001260,
      DO(11) => blk00000001_blk0000092c_sig00001261,
      DO(10) => blk00000001_blk0000092c_sig00001262,
      DO(9) => blk00000001_blk0000092c_sig00001263,
      DO(8) => blk00000001_blk0000092c_sig00001264,
      DO(7) => blk00000001_blk0000092c_sig00001255,
      DO(6) => blk00000001_blk0000092c_sig00001256,
      DO(5) => blk00000001_blk0000092c_sig00001257,
      DO(4) => blk00000001_blk0000092c_sig00001258,
      DO(3) => blk00000001_blk0000092c_sig00001259,
      DO(2) => blk00000001_blk0000092c_sig0000125a,
      DO(1) => blk00000001_blk0000092c_sig0000125b,
      DO(0) => blk00000001_blk0000092c_sig0000125c,
      WRADDR(8) => blk00000001_sig000001d0,
      WRADDR(7) => blk00000001_sig000001cf,
      WRADDR(6) => blk00000001_sig000001ce,
      WRADDR(5) => blk00000001_sig000001cd,
      WRADDR(4) => blk00000001_blk0000092c_sig00001295,
      WRADDR(3) => blk00000001_blk0000092c_sig00001295,
      WRADDR(2) => blk00000001_blk0000092c_sig00001295,
      WRADDR(1) => blk00000001_blk0000092c_sig00001295,
      WRADDR(0) => blk00000001_blk0000092c_sig00001295,
      RDADDR(8) => blk00000001_sig000001c0,
      RDADDR(7) => blk00000001_sig000001bf,
      RDADDR(6) => blk00000001_sig000001be,
      RDADDR(5) => blk00000001_sig000001b9,
      RDADDR(4) => blk00000001_blk0000092c_sig00001295,
      RDADDR(3) => blk00000001_blk0000092c_sig00001295,
      RDADDR(2) => blk00000001_blk0000092c_sig00001295,
      RDADDR(1) => blk00000001_blk0000092c_sig00001295,
      RDADDR(0) => blk00000001_blk0000092c_sig00001295,
      DI(31) => blk00000001_blk0000092c_sig00001295,
      DI(30) => blk00000001_blk0000092c_sig00001295,
      DI(29) => blk00000001_blk0000092c_sig00001295,
      DI(28) => blk00000001_sig000002c0,
      DI(27) => blk00000001_sig000002bf,
      DI(26) => blk00000001_sig000002be,
      DI(25) => blk00000001_sig000002bd,
      DI(24) => blk00000001_sig000002bc,
      DI(23) => blk00000001_sig000002ba,
      DI(22) => blk00000001_sig000002b9,
      DI(21) => blk00000001_sig000002b8,
      DI(20) => blk00000001_sig000002b7,
      DI(19) => blk00000001_sig000002b6,
      DI(18) => blk00000001_sig000002b5,
      DI(17) => blk00000001_sig000002b4,
      DI(16) => blk00000001_sig000002b3,
      DI(15) => blk00000001_sig000002b1,
      DI(14) => blk00000001_sig000002b0,
      DI(13) => blk00000001_sig000002af,
      DI(12) => blk00000001_sig000002ae,
      DI(11) => blk00000001_sig000002ad,
      DI(10) => blk00000001_sig000002ac,
      DI(9) => blk00000001_sig000002ab,
      DI(8) => blk00000001_sig000002aa,
      DI(7) => blk00000001_sig000002a8,
      DI(6) => blk00000001_sig000002a7,
      DI(5) => blk00000001_sig000002a6,
      DI(4) => blk00000001_sig000002a5,
      DI(3) => blk00000001_sig000002a4,
      DI(2) => blk00000001_sig000002a3,
      DI(1) => blk00000001_sig000002a2,
      DI(0) => blk00000001_sig000002a1
    );
  blk00000001_blk0000092c_blk0000094d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126d,
      Q => blk00000001_sig00000240
    );
  blk00000001_blk0000092c_blk0000094c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126e,
      Q => blk00000001_sig0000023f
    );
  blk00000001_blk0000092c_blk0000094b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126f,
      Q => blk00000001_sig0000023e
    );
  blk00000001_blk0000092c_blk0000094a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001270,
      Q => blk00000001_sig0000023d
    );
  blk00000001_blk0000092c_blk00000949 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001271,
      Q => blk00000001_sig0000023c
    );
  blk00000001_blk0000092c_blk00000948 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001274,
      Q => blk00000001_sig0000023b
    );
  blk00000001_blk0000092c_blk00000947 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001265,
      Q => blk00000001_sig0000023a
    );
  blk00000001_blk0000092c_blk00000946 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001266,
      Q => blk00000001_sig00000239
    );
  blk00000001_blk0000092c_blk00000945 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001267,
      Q => blk00000001_sig00000238
    );
  blk00000001_blk0000092c_blk00000944 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001268,
      Q => blk00000001_sig00000237
    );
  blk00000001_blk0000092c_blk00000943 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001269,
      Q => blk00000001_sig00000236
    );
  blk00000001_blk0000092c_blk00000942 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126a,
      Q => blk00000001_sig00000235
    );
  blk00000001_blk0000092c_blk00000941 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126b,
      Q => blk00000001_sig00000234
    );
  blk00000001_blk0000092c_blk00000940 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000126c,
      Q => blk00000001_sig00000233
    );
  blk00000001_blk0000092c_blk0000093f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001273,
      Q => blk00000001_sig00000232
    );
  blk00000001_blk0000092c_blk0000093e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125d,
      Q => blk00000001_sig00000231
    );
  blk00000001_blk0000092c_blk0000093d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125e,
      Q => blk00000001_sig00000230
    );
  blk00000001_blk0000092c_blk0000093c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125f,
      Q => blk00000001_sig0000022f
    );
  blk00000001_blk0000092c_blk0000093b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001260,
      Q => blk00000001_sig0000022e
    );
  blk00000001_blk0000092c_blk0000093a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001261,
      Q => blk00000001_sig0000022d
    );
  blk00000001_blk0000092c_blk00000939 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001262,
      Q => blk00000001_sig0000022c
    );
  blk00000001_blk0000092c_blk00000938 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001263,
      Q => blk00000001_sig0000022b
    );
  blk00000001_blk0000092c_blk00000937 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001264,
      Q => blk00000001_sig0000022a
    );
  blk00000001_blk0000092c_blk00000936 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001272,
      Q => blk00000001_sig00000229
    );
  blk00000001_blk0000092c_blk00000935 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001255,
      Q => blk00000001_sig00000228
    );
  blk00000001_blk0000092c_blk00000934 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001256,
      Q => blk00000001_sig00000227
    );
  blk00000001_blk0000092c_blk00000933 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001257,
      Q => blk00000001_sig00000226
    );
  blk00000001_blk0000092c_blk00000932 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001258,
      Q => blk00000001_sig00000225
    );
  blk00000001_blk0000092c_blk00000931 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig00001259,
      Q => blk00000001_sig00000224
    );
  blk00000001_blk0000092c_blk00000930 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125a,
      Q => blk00000001_sig00000223
    );
  blk00000001_blk0000092c_blk0000092f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125b,
      Q => blk00000001_sig00000222
    );
  blk00000001_blk0000092c_blk0000092e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000092c_sig0000125c,
      Q => blk00000001_sig00000221
    );
  blk00000001_blk0000092c_blk0000092d : GND
    port map (
      G => blk00000001_blk0000092c_sig00001295
    );
  blk00000001_blk0000094f_blk00000971 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000008e,
      RDCLK => aclk,
      WREN => blk00000001_sig0000008e,
      RDEN => blk00000001_sig0000008e,
      WRCLK => aclk,
      SSR => blk00000001_blk0000094f_sig00001302,
      DIP(3) => blk00000001_blk0000094f_sig00001302,
      DIP(2) => blk00000001_sig000002db,
      DIP(1) => blk00000001_sig000002d2,
      DIP(0) => blk00000001_sig000002c9,
      DOP(3) => NLW_blk00000001_blk0000094f_blk00000971_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk0000094f_sig000012e1,
      DOP(1) => blk00000001_blk0000094f_sig000012e0,
      DOP(0) => blk00000001_blk0000094f_sig000012df,
      WE(3) => blk00000001_sig000001d8,
      WE(2) => blk00000001_sig000001d8,
      WE(1) => blk00000001_sig000001d8,
      WE(0) => blk00000001_sig000001d8,
      DO(31) => NLW_blk00000001_blk0000094f_blk00000971_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk0000094f_blk00000971_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk0000094f_blk00000971_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk0000094f_sig000012da,
      DO(27) => blk00000001_blk0000094f_sig000012db,
      DO(26) => blk00000001_blk0000094f_sig000012dc,
      DO(25) => blk00000001_blk0000094f_sig000012dd,
      DO(24) => blk00000001_blk0000094f_sig000012de,
      DO(23) => blk00000001_blk0000094f_sig000012d2,
      DO(22) => blk00000001_blk0000094f_sig000012d3,
      DO(21) => blk00000001_blk0000094f_sig000012d4,
      DO(20) => blk00000001_blk0000094f_sig000012d5,
      DO(19) => blk00000001_blk0000094f_sig000012d6,
      DO(18) => blk00000001_blk0000094f_sig000012d7,
      DO(17) => blk00000001_blk0000094f_sig000012d8,
      DO(16) => blk00000001_blk0000094f_sig000012d9,
      DO(15) => blk00000001_blk0000094f_sig000012ca,
      DO(14) => blk00000001_blk0000094f_sig000012cb,
      DO(13) => blk00000001_blk0000094f_sig000012cc,
      DO(12) => blk00000001_blk0000094f_sig000012cd,
      DO(11) => blk00000001_blk0000094f_sig000012ce,
      DO(10) => blk00000001_blk0000094f_sig000012cf,
      DO(9) => blk00000001_blk0000094f_sig000012d0,
      DO(8) => blk00000001_blk0000094f_sig000012d1,
      DO(7) => blk00000001_blk0000094f_sig000012c2,
      DO(6) => blk00000001_blk0000094f_sig000012c3,
      DO(5) => blk00000001_blk0000094f_sig000012c4,
      DO(4) => blk00000001_blk0000094f_sig000012c5,
      DO(3) => blk00000001_blk0000094f_sig000012c6,
      DO(2) => blk00000001_blk0000094f_sig000012c7,
      DO(1) => blk00000001_blk0000094f_sig000012c8,
      DO(0) => blk00000001_blk0000094f_sig000012c9,
      WRADDR(8) => blk00000001_sig000001d4,
      WRADDR(7) => blk00000001_sig000001d3,
      WRADDR(6) => blk00000001_sig000001d2,
      WRADDR(5) => blk00000001_sig000001d1,
      WRADDR(4) => blk00000001_blk0000094f_sig00001302,
      WRADDR(3) => blk00000001_blk0000094f_sig00001302,
      WRADDR(2) => blk00000001_blk0000094f_sig00001302,
      WRADDR(1) => blk00000001_blk0000094f_sig00001302,
      WRADDR(0) => blk00000001_blk0000094f_sig00001302,
      RDADDR(8) => blk00000001_sig000001c4,
      RDADDR(7) => blk00000001_sig000001c3,
      RDADDR(6) => blk00000001_sig000001c2,
      RDADDR(5) => blk00000001_sig000001c1,
      RDADDR(4) => blk00000001_blk0000094f_sig00001302,
      RDADDR(3) => blk00000001_blk0000094f_sig00001302,
      RDADDR(2) => blk00000001_blk0000094f_sig00001302,
      RDADDR(1) => blk00000001_blk0000094f_sig00001302,
      RDADDR(0) => blk00000001_blk0000094f_sig00001302,
      DI(31) => blk00000001_blk0000094f_sig00001302,
      DI(30) => blk00000001_blk0000094f_sig00001302,
      DI(29) => blk00000001_blk0000094f_sig00001302,
      DI(28) => blk00000001_sig000002e0,
      DI(27) => blk00000001_sig000002df,
      DI(26) => blk00000001_sig000002de,
      DI(25) => blk00000001_sig000002dd,
      DI(24) => blk00000001_sig000002dc,
      DI(23) => blk00000001_sig000002da,
      DI(22) => blk00000001_sig000002d9,
      DI(21) => blk00000001_sig000002d8,
      DI(20) => blk00000001_sig000002d7,
      DI(19) => blk00000001_sig000002d6,
      DI(18) => blk00000001_sig000002d5,
      DI(17) => blk00000001_sig000002d4,
      DI(16) => blk00000001_sig000002d3,
      DI(15) => blk00000001_sig000002d1,
      DI(14) => blk00000001_sig000002d0,
      DI(13) => blk00000001_sig000002cf,
      DI(12) => blk00000001_sig000002ce,
      DI(11) => blk00000001_sig000002cd,
      DI(10) => blk00000001_sig000002cc,
      DI(9) => blk00000001_sig000002cb,
      DI(8) => blk00000001_sig000002ca,
      DI(7) => blk00000001_sig000002c8,
      DI(6) => blk00000001_sig000002c7,
      DI(5) => blk00000001_sig000002c6,
      DI(4) => blk00000001_sig000002c5,
      DI(3) => blk00000001_sig000002c4,
      DI(2) => blk00000001_sig000002c3,
      DI(1) => blk00000001_sig000002c2,
      DI(0) => blk00000001_sig000002c1
    );
  blk00000001_blk0000094f_blk00000970 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012da,
      Q => blk00000001_sig00000260
    );
  blk00000001_blk0000094f_blk0000096f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012db,
      Q => blk00000001_sig0000025f
    );
  blk00000001_blk0000094f_blk0000096e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012dc,
      Q => blk00000001_sig0000025e
    );
  blk00000001_blk0000094f_blk0000096d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012dd,
      Q => blk00000001_sig0000025d
    );
  blk00000001_blk0000094f_blk0000096c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012de,
      Q => blk00000001_sig0000025c
    );
  blk00000001_blk0000094f_blk0000096b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012e1,
      Q => blk00000001_sig0000025b
    );
  blk00000001_blk0000094f_blk0000096a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d2,
      Q => blk00000001_sig0000025a
    );
  blk00000001_blk0000094f_blk00000969 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d3,
      Q => blk00000001_sig00000259
    );
  blk00000001_blk0000094f_blk00000968 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d4,
      Q => blk00000001_sig00000258
    );
  blk00000001_blk0000094f_blk00000967 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d5,
      Q => blk00000001_sig00000257
    );
  blk00000001_blk0000094f_blk00000966 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d6,
      Q => blk00000001_sig00000256
    );
  blk00000001_blk0000094f_blk00000965 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d7,
      Q => blk00000001_sig00000255
    );
  blk00000001_blk0000094f_blk00000964 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d8,
      Q => blk00000001_sig00000254
    );
  blk00000001_blk0000094f_blk00000963 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d9,
      Q => blk00000001_sig00000253
    );
  blk00000001_blk0000094f_blk00000962 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012e0,
      Q => blk00000001_sig00000252
    );
  blk00000001_blk0000094f_blk00000961 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012ca,
      Q => blk00000001_sig00000251
    );
  blk00000001_blk0000094f_blk00000960 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012cb,
      Q => blk00000001_sig00000250
    );
  blk00000001_blk0000094f_blk0000095f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012cc,
      Q => blk00000001_sig0000024f
    );
  blk00000001_blk0000094f_blk0000095e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012cd,
      Q => blk00000001_sig0000024e
    );
  blk00000001_blk0000094f_blk0000095d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012ce,
      Q => blk00000001_sig0000024d
    );
  blk00000001_blk0000094f_blk0000095c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012cf,
      Q => blk00000001_sig0000024c
    );
  blk00000001_blk0000094f_blk0000095b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d0,
      Q => blk00000001_sig0000024b
    );
  blk00000001_blk0000094f_blk0000095a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012d1,
      Q => blk00000001_sig0000024a
    );
  blk00000001_blk0000094f_blk00000959 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012df,
      Q => blk00000001_sig00000249
    );
  blk00000001_blk0000094f_blk00000958 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c2,
      Q => blk00000001_sig00000248
    );
  blk00000001_blk0000094f_blk00000957 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c3,
      Q => blk00000001_sig00000247
    );
  blk00000001_blk0000094f_blk00000956 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c4,
      Q => blk00000001_sig00000246
    );
  blk00000001_blk0000094f_blk00000955 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c5,
      Q => blk00000001_sig00000245
    );
  blk00000001_blk0000094f_blk00000954 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c6,
      Q => blk00000001_sig00000244
    );
  blk00000001_blk0000094f_blk00000953 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c7,
      Q => blk00000001_sig00000243
    );
  blk00000001_blk0000094f_blk00000952 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c8,
      Q => blk00000001_sig00000242
    );
  blk00000001_blk0000094f_blk00000951 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000094f_sig000012c9,
      Q => blk00000001_sig00000241
    );
  blk00000001_blk0000094f_blk00000950 : GND
    port map (
      G => blk00000001_blk0000094f_sig00001302
    );
  blk00000001_blk00000972_blk00000973_blk00000977 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000972_blk00000973_sig0000130e,
      Q => blk00000001_sig00000da6
    );
  blk00000001_blk00000972_blk00000973_blk00000976 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000972_blk00000973_sig0000130d,
      A1 => blk00000001_blk00000972_blk00000973_sig0000130c,
      A2 => blk00000001_blk00000972_blk00000973_sig0000130c,
      A3 => blk00000001_blk00000972_blk00000973_sig0000130c,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000001a6,
      Q => blk00000001_blk00000972_blk00000973_sig0000130e,
      Q15 => NLW_blk00000001_blk00000972_blk00000973_blk00000976_Q15_UNCONNECTED
    );
  blk00000001_blk00000972_blk00000973_blk00000975 : VCC
    port map (
      P => blk00000001_blk00000972_blk00000973_sig0000130d
    );
  blk00000001_blk00000972_blk00000973_blk00000974 : GND
    port map (
      G => blk00000001_blk00000972_blk00000973_sig0000130c
    );
  blk00000001_blk00000978_blk00000979_blk0000097d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000978_blk00000979_sig0000131a,
      Q => blk00000001_sig00000ddc
    );
  blk00000001_blk00000978_blk00000979_blk0000097c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000978_blk00000979_sig00001319,
      A1 => blk00000001_blk00000978_blk00000979_sig00001318,
      A2 => blk00000001_blk00000978_blk00000979_sig00001318,
      A3 => blk00000001_blk00000978_blk00000979_sig00001318,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000ddd,
      Q => blk00000001_blk00000978_blk00000979_sig0000131a,
      Q15 => NLW_blk00000001_blk00000978_blk00000979_blk0000097c_Q15_UNCONNECTED
    );
  blk00000001_blk00000978_blk00000979_blk0000097b : VCC
    port map (
      P => blk00000001_blk00000978_blk00000979_sig00001319
    );
  blk00000001_blk00000978_blk00000979_blk0000097a : GND
    port map (
      G => blk00000001_blk00000978_blk00000979_sig00001318
    );
  blk00000001_blk0000097e_blk0000097f_blk00000983 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000097e_blk0000097f_sig00001326,
      Q => blk00000001_sig00000dde
    );
  blk00000001_blk0000097e_blk0000097f_blk00000982 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000097e_blk0000097f_sig00001325,
      A1 => blk00000001_blk0000097e_blk0000097f_sig00001324,
      A2 => blk00000001_blk0000097e_blk0000097f_sig00001324,
      A3 => blk00000001_blk0000097e_blk0000097f_sig00001324,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dec,
      Q => blk00000001_blk0000097e_blk0000097f_sig00001326,
      Q15 => NLW_blk00000001_blk0000097e_blk0000097f_blk00000982_Q15_UNCONNECTED
    );
  blk00000001_blk0000097e_blk0000097f_blk00000981 : VCC
    port map (
      P => blk00000001_blk0000097e_blk0000097f_sig00001325
    );
  blk00000001_blk0000097e_blk0000097f_blk00000980 : GND
    port map (
      G => blk00000001_blk0000097e_blk0000097f_sig00001324
    );
  blk00000001_blk00000984_blk00000985_blk00000989 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000984_blk00000985_sig00001332,
      Q => blk00000001_sig00000de7
    );
  blk00000001_blk00000984_blk00000985_blk00000988 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000984_blk00000985_sig00001331,
      A1 => blk00000001_blk00000984_blk00000985_sig00001330,
      A2 => blk00000001_blk00000984_blk00000985_sig00001330,
      A3 => blk00000001_blk00000984_blk00000985_sig00001330,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000000bb,
      Q => blk00000001_blk00000984_blk00000985_sig00001332,
      Q15 => NLW_blk00000001_blk00000984_blk00000985_blk00000988_Q15_UNCONNECTED
    );
  blk00000001_blk00000984_blk00000985_blk00000987 : VCC
    port map (
      P => blk00000001_blk00000984_blk00000985_sig00001331
    );
  blk00000001_blk00000984_blk00000985_blk00000986 : GND
    port map (
      G => blk00000001_blk00000984_blk00000985_sig00001330
    );
  blk00000001_blk0000098a_blk0000098b_blk0000098f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk0000098a_blk0000098b_sig0000133e,
      Q => blk00000001_sig000001af
    );
  blk00000001_blk0000098a_blk0000098b_blk0000098e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk0000098a_blk0000098b_sig0000133d,
      A1 => blk00000001_blk0000098a_blk0000098b_sig0000133c,
      A2 => blk00000001_blk0000098a_blk0000098b_sig0000133c,
      A3 => blk00000001_blk0000098a_blk0000098b_sig0000133c,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000000bb,
      Q => blk00000001_blk0000098a_blk0000098b_sig0000133e,
      Q15 => NLW_blk00000001_blk0000098a_blk0000098b_blk0000098e_Q15_UNCONNECTED
    );
  blk00000001_blk0000098a_blk0000098b_blk0000098d : VCC
    port map (
      P => blk00000001_blk0000098a_blk0000098b_sig0000133d
    );
  blk00000001_blk0000098a_blk0000098b_blk0000098c : GND
    port map (
      G => blk00000001_blk0000098a_blk0000098b_sig0000133c
    );
  blk00000001_blk000009c5_blk000009d7 : INV
    port map (
      I => blk00000001_sig00000e3c,
      O => blk00000001_blk000009c5_sig00001352
    );
  blk00000001_blk000009c5_blk000009d6 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e3d,
      O => blk00000001_blk000009c5_sig00001356
    );
  blk00000001_blk000009c5_blk000009d5 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e3e,
      O => blk00000001_blk000009c5_sig00001355
    );
  blk00000001_blk000009c5_blk000009d4 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e3f,
      O => blk00000001_blk000009c5_sig00001354
    );
  blk00000001_blk000009c5_blk000009d3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e40,
      O => blk00000001_blk000009c5_sig00001353
    );
  blk00000001_blk000009c5_blk000009d2 : MUXCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134c,
      DI => blk00000001_blk000009c5_sig0000134b,
      S => blk00000001_blk000009c5_sig00001352,
      O => blk00000001_blk000009c5_sig00001351
    );
  blk00000001_blk000009c5_blk000009d1 : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134c,
      LI => blk00000001_blk000009c5_sig00001352,
      O => blk00000001_sig00000e35
    );
  blk00000001_blk000009c5_blk000009d0 : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134d,
      LI => blk00000001_sig00000e41,
      O => blk00000001_sig00000e3a
    );
  blk00000001_blk000009c5_blk000009cf : MUXCY
    port map (
      CI => blk00000001_blk000009c5_sig00001351,
      DI => blk00000001_blk000009c5_sig0000134c,
      S => blk00000001_blk000009c5_sig00001356,
      O => blk00000001_blk000009c5_sig00001350
    );
  blk00000001_blk000009c5_blk000009ce : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig00001351,
      LI => blk00000001_blk000009c5_sig00001356,
      O => blk00000001_sig00000e36
    );
  blk00000001_blk000009c5_blk000009cd : MUXCY
    port map (
      CI => blk00000001_blk000009c5_sig00001350,
      DI => blk00000001_blk000009c5_sig0000134c,
      S => blk00000001_blk000009c5_sig00001355,
      O => blk00000001_blk000009c5_sig0000134f
    );
  blk00000001_blk000009c5_blk000009cc : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig00001350,
      LI => blk00000001_blk000009c5_sig00001355,
      O => blk00000001_sig00000e37
    );
  blk00000001_blk000009c5_blk000009cb : MUXCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134f,
      DI => blk00000001_blk000009c5_sig0000134c,
      S => blk00000001_blk000009c5_sig00001354,
      O => blk00000001_blk000009c5_sig0000134e
    );
  blk00000001_blk000009c5_blk000009ca : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134f,
      LI => blk00000001_blk000009c5_sig00001354,
      O => blk00000001_sig00000e38
    );
  blk00000001_blk000009c5_blk000009c9 : MUXCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134e,
      DI => blk00000001_blk000009c5_sig0000134c,
      S => blk00000001_blk000009c5_sig00001353,
      O => blk00000001_blk000009c5_sig0000134d
    );
  blk00000001_blk000009c5_blk000009c8 : XORCY
    port map (
      CI => blk00000001_blk000009c5_sig0000134e,
      LI => blk00000001_blk000009c5_sig00001353,
      O => blk00000001_sig00000e39
    );
  blk00000001_blk000009c5_blk000009c7 : GND
    port map (
      G => blk00000001_blk000009c5_sig0000134c
    );
  blk00000001_blk000009c5_blk000009c6 : VCC
    port map (
      P => blk00000001_blk000009c5_sig0000134b
    );
  blk00000001_blk000009e2_blk000009ee : INV
    port map (
      I => blk00000001_sig00000e4b,
      O => blk00000001_blk000009e2_sig00001364
    );
  blk00000001_blk000009e2_blk000009ed : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e4c,
      O => blk00000001_blk000009e2_sig00001366
    );
  blk00000001_blk000009e2_blk000009ec : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e4d,
      O => blk00000001_blk000009e2_sig00001365
    );
  blk00000001_blk000009e2_blk000009eb : MUXCY
    port map (
      CI => blk00000001_blk000009e2_sig00001360,
      DI => blk00000001_blk000009e2_sig0000135f,
      S => blk00000001_blk000009e2_sig00001364,
      O => blk00000001_blk000009e2_sig00001363
    );
  blk00000001_blk000009e2_blk000009ea : XORCY
    port map (
      CI => blk00000001_blk000009e2_sig00001360,
      LI => blk00000001_blk000009e2_sig00001364,
      O => blk00000001_sig00000e46
    );
  blk00000001_blk000009e2_blk000009e9 : XORCY
    port map (
      CI => blk00000001_blk000009e2_sig00001361,
      LI => blk00000001_sig00000e4e,
      O => blk00000001_sig00000e49
    );
  blk00000001_blk000009e2_blk000009e8 : MUXCY
    port map (
      CI => blk00000001_blk000009e2_sig00001363,
      DI => blk00000001_blk000009e2_sig00001360,
      S => blk00000001_blk000009e2_sig00001366,
      O => blk00000001_blk000009e2_sig00001362
    );
  blk00000001_blk000009e2_blk000009e7 : XORCY
    port map (
      CI => blk00000001_blk000009e2_sig00001363,
      LI => blk00000001_blk000009e2_sig00001366,
      O => blk00000001_sig00000e47
    );
  blk00000001_blk000009e2_blk000009e6 : MUXCY
    port map (
      CI => blk00000001_blk000009e2_sig00001362,
      DI => blk00000001_blk000009e2_sig00001360,
      S => blk00000001_blk000009e2_sig00001365,
      O => blk00000001_blk000009e2_sig00001361
    );
  blk00000001_blk000009e2_blk000009e5 : XORCY
    port map (
      CI => blk00000001_blk000009e2_sig00001362,
      LI => blk00000001_blk000009e2_sig00001365,
      O => blk00000001_sig00000e48
    );
  blk00000001_blk000009e2_blk000009e4 : GND
    port map (
      G => blk00000001_blk000009e2_sig00001360
    );
  blk00000001_blk000009e2_blk000009e3 : VCC
    port map (
      P => blk00000001_blk000009e2_sig0000135f
    );
  blk00000001_blk000009fb_blk00000a0a : INV
    port map (
      I => blk00000001_sig00000e59,
      O => blk00000001_blk000009fb_sig00001377
    );
  blk00000001_blk000009fb_blk00000a09 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e5a,
      O => blk00000001_blk000009fb_sig0000137a
    );
  blk00000001_blk000009fb_blk00000a08 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e5b,
      O => blk00000001_blk000009fb_sig00001379
    );
  blk00000001_blk000009fb_blk00000a07 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e5c,
      O => blk00000001_blk000009fb_sig00001378
    );
  blk00000001_blk000009fb_blk00000a06 : MUXCY
    port map (
      CI => blk00000001_blk000009fb_sig00001372,
      DI => blk00000001_blk000009fb_sig00001371,
      S => blk00000001_blk000009fb_sig00001377,
      O => blk00000001_blk000009fb_sig00001376
    );
  blk00000001_blk000009fb_blk00000a05 : XORCY
    port map (
      CI => blk00000001_blk000009fb_sig00001372,
      LI => blk00000001_blk000009fb_sig00001377,
      O => blk00000001_sig00000e53
    );
  blk00000001_blk000009fb_blk00000a04 : XORCY
    port map (
      CI => blk00000001_blk000009fb_sig00001373,
      LI => blk00000001_sig00000e5d,
      O => blk00000001_sig00000e57
    );
  blk00000001_blk000009fb_blk00000a03 : MUXCY
    port map (
      CI => blk00000001_blk000009fb_sig00001376,
      DI => blk00000001_blk000009fb_sig00001372,
      S => blk00000001_blk000009fb_sig0000137a,
      O => blk00000001_blk000009fb_sig00001375
    );
  blk00000001_blk000009fb_blk00000a02 : XORCY
    port map (
      CI => blk00000001_blk000009fb_sig00001376,
      LI => blk00000001_blk000009fb_sig0000137a,
      O => blk00000001_sig00000e54
    );
  blk00000001_blk000009fb_blk00000a01 : MUXCY
    port map (
      CI => blk00000001_blk000009fb_sig00001375,
      DI => blk00000001_blk000009fb_sig00001372,
      S => blk00000001_blk000009fb_sig00001379,
      O => blk00000001_blk000009fb_sig00001374
    );
  blk00000001_blk000009fb_blk00000a00 : XORCY
    port map (
      CI => blk00000001_blk000009fb_sig00001375,
      LI => blk00000001_blk000009fb_sig00001379,
      O => blk00000001_sig00000e55
    );
  blk00000001_blk000009fb_blk000009ff : MUXCY
    port map (
      CI => blk00000001_blk000009fb_sig00001374,
      DI => blk00000001_blk000009fb_sig00001372,
      S => blk00000001_blk000009fb_sig00001378,
      O => blk00000001_blk000009fb_sig00001373
    );
  blk00000001_blk000009fb_blk000009fe : XORCY
    port map (
      CI => blk00000001_blk000009fb_sig00001374,
      LI => blk00000001_blk000009fb_sig00001378,
      O => blk00000001_sig00000e56
    );
  blk00000001_blk000009fb_blk000009fd : GND
    port map (
      G => blk00000001_blk000009fb_sig00001372
    );
  blk00000001_blk000009fb_blk000009fc : VCC
    port map (
      P => blk00000001_blk000009fb_sig00001371
    );
  blk00000001_blk00000a0b_blk00000a0c_blk00000a10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a0b_blk00000a0c_sig00001385,
      Q => blk00000001_sig00000e23
    );
  blk00000001_blk00000a0b_blk00000a0c_blk00000a0f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000a0b_blk00000a0c_sig00001384,
      A1 => blk00000001_blk00000a0b_blk00000a0c_sig00001383,
      A2 => blk00000001_blk00000a0b_blk00000a0c_sig00001384,
      A3 => blk00000001_blk00000a0b_blk00000a0c_sig00001383,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000e1e,
      Q => blk00000001_blk00000a0b_blk00000a0c_sig00001385,
      Q15 => NLW_blk00000001_blk00000a0b_blk00000a0c_blk00000a0f_Q15_UNCONNECTED
    );
  blk00000001_blk00000a0b_blk00000a0c_blk00000a0e : VCC
    port map (
      P => blk00000001_blk00000a0b_blk00000a0c_sig00001384
    );
  blk00000001_blk00000a0b_blk00000a0c_blk00000a0d : GND
    port map (
      G => blk00000001_blk00000a0b_blk00000a0c_sig00001383
    );
  blk00000001_blk00000a15_blk00000a1e : INV
    port map (
      I => blk00000001_sig00000e6a,
      O => blk00000001_blk00000a15_sig00001390
    );
  blk00000001_blk00000a15_blk00000a1d : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000e6b,
      O => blk00000001_blk00000a15_sig00001391
    );
  blk00000001_blk00000a15_blk00000a1c : MUXCY
    port map (
      CI => blk00000001_blk00000a15_sig0000138d,
      DI => blk00000001_blk00000a15_sig0000138c,
      S => blk00000001_blk00000a15_sig00001390,
      O => blk00000001_blk00000a15_sig0000138f
    );
  blk00000001_blk00000a15_blk00000a1b : XORCY
    port map (
      CI => blk00000001_blk00000a15_sig0000138d,
      LI => blk00000001_blk00000a15_sig00001390,
      O => blk00000001_sig00000e67
    );
  blk00000001_blk00000a15_blk00000a1a : XORCY
    port map (
      CI => blk00000001_blk00000a15_sig0000138e,
      LI => blk00000001_sig00000e6c,
      O => blk00000001_sig00000e69
    );
  blk00000001_blk00000a15_blk00000a19 : MUXCY
    port map (
      CI => blk00000001_blk00000a15_sig0000138f,
      DI => blk00000001_blk00000a15_sig0000138d,
      S => blk00000001_blk00000a15_sig00001391,
      O => blk00000001_blk00000a15_sig0000138e
    );
  blk00000001_blk00000a15_blk00000a18 : XORCY
    port map (
      CI => blk00000001_blk00000a15_sig0000138f,
      LI => blk00000001_blk00000a15_sig00001391,
      O => blk00000001_sig00000e68
    );
  blk00000001_blk00000a15_blk00000a17 : GND
    port map (
      G => blk00000001_blk00000a15_sig0000138d
    );
  blk00000001_blk00000a15_blk00000a16 : VCC
    port map (
      P => blk00000001_blk00000a15_sig0000138c
    );
  blk00000001_blk00000a1f_blk00000a20_blk00000a24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a1f_blk00000a20_sig000013a5,
      Q => blk00000001_sig00000e20
    );
  blk00000001_blk00000a1f_blk00000a20_blk00000a23 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000e21,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000a1f_blk00000a20_sig000013a5,
      Q31 => NLW_blk00000001_blk00000a1f_blk00000a20_blk00000a23_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000a1f_blk00000a20_sig000013a4,
      A(3) => blk00000001_blk00000a1f_blk00000a20_sig000013a3,
      A(2) => blk00000001_blk00000a1f_blk00000a20_sig000013a4,
      A(1) => blk00000001_blk00000a1f_blk00000a20_sig000013a3,
      A(0) => blk00000001_blk00000a1f_blk00000a20_sig000013a3
    );
  blk00000001_blk00000a1f_blk00000a20_blk00000a22 : VCC
    port map (
      P => blk00000001_blk00000a1f_blk00000a20_sig000013a4
    );
  blk00000001_blk00000a1f_blk00000a20_blk00000a21 : GND
    port map (
      G => blk00000001_blk00000a1f_blk00000a20_sig000013a3
    );
  blk00000001_blk00000a25_blk00000a26_blk00000a2a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a25_blk00000a26_sig000013b0,
      Q => blk00000001_sig00000de8
    );
  blk00000001_blk00000a25_blk00000a26_blk00000a29 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000a25_blk00000a26_sig000013ae,
      A1 => blk00000001_blk00000a25_blk00000a26_sig000013ae,
      A2 => blk00000001_blk00000a25_blk00000a26_sig000013af,
      A3 => blk00000001_blk00000a25_blk00000a26_sig000013ae,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dec,
      Q => blk00000001_blk00000a25_blk00000a26_sig000013b0,
      Q15 => NLW_blk00000001_blk00000a25_blk00000a26_blk00000a29_Q15_UNCONNECTED
    );
  blk00000001_blk00000a25_blk00000a26_blk00000a28 : VCC
    port map (
      P => blk00000001_blk00000a25_blk00000a26_sig000013af
    );
  blk00000001_blk00000a25_blk00000a26_blk00000a27 : GND
    port map (
      G => blk00000001_blk00000a25_blk00000a26_sig000013ae
    );
  blk00000001_blk00000a2b_blk00000a2c_blk00000a30 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a2b_blk00000a2c_sig000013bb,
      Q => blk00000001_sig000001ad
    );
  blk00000001_blk00000a2b_blk00000a2c_blk00000a2f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000a2b_blk00000a2c_sig000013ba,
      A1 => blk00000001_blk00000a2b_blk00000a2c_sig000013ba,
      A2 => blk00000001_blk00000a2b_blk00000a2c_sig000013b9,
      A3 => blk00000001_blk00000a2b_blk00000a2c_sig000013ba,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig000000c0,
      Q => blk00000001_blk00000a2b_blk00000a2c_sig000013bb,
      Q15 => NLW_blk00000001_blk00000a2b_blk00000a2c_blk00000a2f_Q15_UNCONNECTED
    );
  blk00000001_blk00000a2b_blk00000a2c_blk00000a2e : VCC
    port map (
      P => blk00000001_blk00000a2b_blk00000a2c_sig000013ba
    );
  blk00000001_blk00000a2b_blk00000a2c_blk00000a2d : GND
    port map (
      G => blk00000001_blk00000a2b_blk00000a2c_sig000013b9
    );
  blk00000001_blk00000a31_blk00000a32_blk00000a36 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a31_blk00000a32_sig000013c6,
      Q => blk00000001_sig000001ac
    );
  blk00000001_blk00000a31_blk00000a32_blk00000a35 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig000000c0,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000a31_blk00000a32_sig000013c6,
      Q31 => NLW_blk00000001_blk00000a31_blk00000a32_blk00000a35_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000a31_blk00000a32_sig000013c5,
      A(3) => blk00000001_blk00000a31_blk00000a32_sig000013c4,
      A(2) => blk00000001_blk00000a31_blk00000a32_sig000013c4,
      A(1) => blk00000001_blk00000a31_blk00000a32_sig000013c5,
      A(0) => blk00000001_blk00000a31_blk00000a32_sig000013c4
    );
  blk00000001_blk00000a31_blk00000a32_blk00000a34 : VCC
    port map (
      P => blk00000001_blk00000a31_blk00000a32_sig000013c5
    );
  blk00000001_blk00000a31_blk00000a32_blk00000a33 : GND
    port map (
      G => blk00000001_blk00000a31_blk00000a32_sig000013c4
    );
  blk00000001_blk00000a37_blk00000a38_blk00000a3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a37_blk00000a38_sig000013da,
      Q => blk00000001_sig000001aa
    );
  blk00000001_blk00000a37_blk00000a38_blk00000a3b : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000deb,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000a37_blk00000a38_sig000013da,
      Q31 => NLW_blk00000001_blk00000a37_blk00000a38_blk00000a3b_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000a37_blk00000a38_sig000013d9,
      A(3) => blk00000001_blk00000a37_blk00000a38_sig000013d8,
      A(2) => blk00000001_blk00000a37_blk00000a38_sig000013d9,
      A(1) => blk00000001_blk00000a37_blk00000a38_sig000013d8,
      A(0) => blk00000001_blk00000a37_blk00000a38_sig000013d8
    );
  blk00000001_blk00000a37_blk00000a38_blk00000a3a : VCC
    port map (
      P => blk00000001_blk00000a37_blk00000a38_sig000013d9
    );
  blk00000001_blk00000a37_blk00000a38_blk00000a39 : GND
    port map (
      G => blk00000001_blk00000a37_blk00000a38_sig000013d8
    );
  blk00000001_blk00000a3d_blk00000a3e_blk00000a42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a3d_blk00000a3e_sig000013ee,
      Q => blk00000001_sig000001a9
    );
  blk00000001_blk00000a3d_blk00000a3e_blk00000a41 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000ded,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000a3d_blk00000a3e_sig000013ee,
      Q31 => NLW_blk00000001_blk00000a3d_blk00000a3e_blk00000a41_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000a3d_blk00000a3e_sig000013ed,
      A(3) => blk00000001_blk00000a3d_blk00000a3e_sig000013ec,
      A(2) => blk00000001_blk00000a3d_blk00000a3e_sig000013ed,
      A(1) => blk00000001_blk00000a3d_blk00000a3e_sig000013ec,
      A(0) => blk00000001_blk00000a3d_blk00000a3e_sig000013ec
    );
  blk00000001_blk00000a3d_blk00000a3e_blk00000a40 : VCC
    port map (
      P => blk00000001_blk00000a3d_blk00000a3e_sig000013ed
    );
  blk00000001_blk00000a3d_blk00000a3e_blk00000a3f : GND
    port map (
      G => blk00000001_blk00000a3d_blk00000a3e_sig000013ec
    );
  blk00000001_blk00000a61_blk00000a62_blk00000a66 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000deb,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000a61_blk00000a62_sig000013f9,
      Q31 => NLW_blk00000001_blk00000a61_blk00000a62_blk00000a66_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000a61_blk00000a62_sig000013fb,
      A(3) => blk00000001_blk00000a61_blk00000a62_sig000013fa,
      A(2) => blk00000001_blk00000a61_blk00000a62_sig000013fb,
      A(1) => blk00000001_blk00000a61_blk00000a62_sig000013fa,
      A(0) => blk00000001_blk00000a61_blk00000a62_sig000013fa
    );
  blk00000001_blk00000a61_blk00000a62_blk00000a65 : VCC
    port map (
      P => blk00000001_blk00000a61_blk00000a62_sig000013fb
    );
  blk00000001_blk00000a61_blk00000a62_blk00000a64 : GND
    port map (
      G => blk00000001_blk00000a61_blk00000a62_sig000013fa
    );
  blk00000001_blk00000a61_blk00000a62_blk00000a63 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a61_blk00000a62_sig000013f9,
      R => blk00000001_sig00000de9,
      Q => blk00000001_sig00000de0
    );
  blk00000001_blk00000a67_blk00000a68_blk00000a6c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a67_blk00000a68_sig00001406,
      Q => blk00000001_sig00000ddf
    );
  blk00000001_blk00000a67_blk00000a68_blk00000a6b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000a67_blk00000a68_sig00001404,
      A1 => blk00000001_blk00000a67_blk00000a68_sig00001405,
      A2 => blk00000001_blk00000a67_blk00000a68_sig00001405,
      A3 => blk00000001_blk00000a67_blk00000a68_sig00001404,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000deb,
      Q => blk00000001_blk00000a67_blk00000a68_sig00001406,
      Q15 => NLW_blk00000001_blk00000a67_blk00000a68_blk00000a6b_Q15_UNCONNECTED
    );
  blk00000001_blk00000a67_blk00000a68_blk00000a6a : VCC
    port map (
      P => blk00000001_blk00000a67_blk00000a68_sig00001405
    );
  blk00000001_blk00000a67_blk00000a68_blk00000a69 : GND
    port map (
      G => blk00000001_blk00000a67_blk00000a68_sig00001404
    );
  blk00000001_blk00000a6d_blk00000a6e_blk00000a72 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000a6d_blk00000a6e_sig00001412,
      A1 => blk00000001_blk00000a6d_blk00000a6e_sig00001413,
      A2 => blk00000001_blk00000a6d_blk00000a6e_sig00001413,
      A3 => blk00000001_blk00000a6d_blk00000a6e_sig00001412,
      CE => blk00000001_sig0000008e,
      CLK => aclk,
      D => blk00000001_sig00000dec,
      Q => blk00000001_blk00000a6d_blk00000a6e_sig00001411,
      Q15 => NLW_blk00000001_blk00000a6d_blk00000a6e_blk00000a72_Q15_UNCONNECTED
    );
  blk00000001_blk00000a6d_blk00000a6e_blk00000a71 : VCC
    port map (
      P => blk00000001_blk00000a6d_blk00000a6e_sig00001413
    );
  blk00000001_blk00000a6d_blk00000a6e_blk00000a70 : GND
    port map (
      G => blk00000001_blk00000a6d_blk00000a6e_sig00001412
    );
  blk00000001_blk00000a6d_blk00000a6e_blk00000a6f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a6d_blk00000a6e_sig00001411,
      R => blk00000001_sig000001ab,
      Q => blk00000001_sig000000be
    );
  blk00000001_blk00000a9e_blk00000ab1 : INV
    port map (
      I => blk00000001_sig00000eb2,
      O => blk00000001_blk00000a9e_sig00001428
    );
  blk00000001_blk00000a9e_blk00000ab0 : INV
    port map (
      I => blk00000001_sig00000eb1,
      O => blk00000001_blk00000a9e_sig00001425
    );
  blk00000001_blk00000a9e_blk00000aaf : INV
    port map (
      I => blk00000001_sig00000eb0,
      O => blk00000001_blk00000a9e_sig00001426
    );
  blk00000001_blk00000a9e_blk00000aae : INV
    port map (
      I => blk00000001_sig00000eaf,
      O => blk00000001_blk00000a9e_sig00001427
    );
  blk00000001_blk00000a9e_blk00000aad : INV
    port map (
      I => blk00000001_sig00000eaf,
      O => blk00000001_blk00000a9e_sig00001429
    );
  blk00000001_blk00000a9e_blk00000aac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a9e_sig00001421,
      Q => blk00000001_sig00000ea2
    );
  blk00000001_blk00000a9e_blk00000aab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a9e_sig00001424,
      Q => blk00000001_sig00000ea3
    );
  blk00000001_blk00000a9e_blk00000aaa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a9e_sig00001423,
      Q => blk00000001_sig00000ea4
    );
  blk00000001_blk00000a9e_blk00000aa9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000a9e_sig00001422,
      Q => blk00000001_sig00000ea5
    );
  blk00000001_blk00000a9e_blk00000aa8 : MUXCY
    port map (
      CI => blk00000001_blk00000a9e_sig00001420,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_blk00000a9e_sig00001429,
      O => blk00000001_blk00000a9e_sig0000142d
    );
  blk00000001_blk00000a9e_blk00000aa7 : MUXCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142d,
      DI => blk00000001_sig00000eaf,
      S => blk00000001_blk00000a9e_sig00001427,
      O => blk00000001_blk00000a9e_sig0000142c
    );
  blk00000001_blk00000a9e_blk00000aa6 : MUXCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142c,
      DI => blk00000001_sig00000eb0,
      S => blk00000001_blk00000a9e_sig00001426,
      O => blk00000001_blk00000a9e_sig0000142b
    );
  blk00000001_blk00000a9e_blk00000aa5 : MUXCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142b,
      DI => blk00000001_sig00000eb1,
      S => blk00000001_blk00000a9e_sig00001425,
      O => blk00000001_blk00000a9e_sig0000142a
    );
  blk00000001_blk00000a9e_blk00000aa4 : XORCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142d,
      LI => blk00000001_blk00000a9e_sig00001427,
      O => blk00000001_blk00000a9e_sig00001424
    );
  blk00000001_blk00000a9e_blk00000aa3 : XORCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142c,
      LI => blk00000001_blk00000a9e_sig00001426,
      O => blk00000001_blk00000a9e_sig00001423
    );
  blk00000001_blk00000a9e_blk00000aa2 : XORCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142b,
      LI => blk00000001_blk00000a9e_sig00001425,
      O => blk00000001_blk00000a9e_sig00001422
    );
  blk00000001_blk00000a9e_blk00000aa1 : XORCY
    port map (
      CI => blk00000001_blk00000a9e_sig0000142a,
      LI => blk00000001_blk00000a9e_sig00001428,
      O => NLW_blk00000001_blk00000a9e_blk00000aa1_O_UNCONNECTED
    );
  blk00000001_blk00000a9e_blk00000aa0 : XORCY
    port map (
      CI => blk00000001_blk00000a9e_sig00001420,
      LI => blk00000001_blk00000a9e_sig00001429,
      O => blk00000001_blk00000a9e_sig00001421
    );
  blk00000001_blk00000a9e_blk00000a9f : VCC
    port map (
      P => blk00000001_blk00000a9e_sig00001420
    );
  blk00000001_blk00000b3c_blk00000b4d : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000ef5,
      O => blk00000001_blk00000b3c_sig00001447
    );
  blk00000001_blk00000b3c_blk00000b4c : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig00000ef2,
      O => blk00000001_blk00000b3c_sig00001446
    );
  blk00000001_blk00000b3c_blk00000b4b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ef2,
      I1 => blk00000001_sig00000ef3,
      O => blk00000001_blk00000b3c_sig0000143e
    );
  blk00000001_blk00000b3c_blk00000b4a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ef3,
      I1 => blk00000001_sig00000ef4,
      O => blk00000001_blk00000b3c_sig0000143f
    );
  blk00000001_blk00000b3c_blk00000b49 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_sig00000ef4,
      I1 => blk00000001_sig00000ef5,
      O => blk00000001_blk00000b3c_sig00001440
    );
  blk00000001_blk00000b3c_blk00000b48 : MUXCY
    port map (
      CI => blk00000001_blk00000b3c_sig0000143d,
      DI => blk00000001_sig00000ef5,
      S => blk00000001_blk00000b3c_sig00001447,
      O => blk00000001_blk00000b3c_sig00001445
    );
  blk00000001_blk00000b3c_blk00000b47 : MUXCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001445,
      DI => blk00000001_sig00000ef4,
      S => blk00000001_blk00000b3c_sig00001440,
      O => blk00000001_blk00000b3c_sig00001444
    );
  blk00000001_blk00000b3c_blk00000b46 : MUXCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001444,
      DI => blk00000001_sig00000ef3,
      S => blk00000001_blk00000b3c_sig0000143f,
      O => blk00000001_blk00000b3c_sig00001443
    );
  blk00000001_blk00000b3c_blk00000b45 : MUXCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001443,
      DI => blk00000001_sig00000ef2,
      S => blk00000001_blk00000b3c_sig0000143e,
      O => blk00000001_blk00000b3c_sig00001442
    );
  blk00000001_blk00000b3c_blk00000b44 : MUXCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001442,
      DI => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_blk00000b3c_sig00001446,
      O => blk00000001_blk00000b3c_sig00001441
    );
  blk00000001_blk00000b3c_blk00000b43 : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001445,
      LI => blk00000001_blk00000b3c_sig00001440,
      O => blk00000001_sig00000ef7
    );
  blk00000001_blk00000b3c_blk00000b42 : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001444,
      LI => blk00000001_blk00000b3c_sig0000143f,
      O => blk00000001_sig00000ef8
    );
  blk00000001_blk00000b3c_blk00000b41 : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001443,
      LI => blk00000001_blk00000b3c_sig0000143e,
      O => blk00000001_sig00000ef9
    );
  blk00000001_blk00000b3c_blk00000b40 : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001442,
      LI => blk00000001_blk00000b3c_sig00001446,
      O => blk00000001_sig00000efa
    );
  blk00000001_blk00000b3c_blk00000b3f : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig00001441,
      LI => blk00000001_blk00000b3c_sig0000143d,
      O => blk00000001_sig00000efb
    );
  blk00000001_blk00000b3c_blk00000b3e : XORCY
    port map (
      CI => blk00000001_blk00000b3c_sig0000143d,
      LI => blk00000001_blk00000b3c_sig00001447,
      O => blk00000001_sig00000ef6
    );
  blk00000001_blk00000b3c_blk00000b3d : GND
    port map (
      G => blk00000001_blk00000b3c_sig0000143d
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b59 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b4e_blk00000b4f_sig00001462,
      Q => blk00000001_sig00000db6
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b58 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd3,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b4e_blk00000b4f_sig00001462,
      Q31 => NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b58_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b4e_blk00000b4f_sig0000145e,
      A(3) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(2) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(1) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(0) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b57 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b4e_blk00000b4f_sig00001461,
      Q => blk00000001_sig00000db5
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b56 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd2,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b4e_blk00000b4f_sig00001461,
      Q31 => NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b56_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b4e_blk00000b4f_sig0000145e,
      A(3) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(2) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(1) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(0) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b55 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b4e_blk00000b4f_sig00001460,
      Q => blk00000001_sig00000db4
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b54 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd1,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b4e_blk00000b4f_sig00001460,
      Q31 => NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b54_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b4e_blk00000b4f_sig0000145e,
      A(3) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(2) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(1) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(0) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b53 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b4e_blk00000b4f_sig0000145f,
      Q => blk00000001_sig00000db3
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b52 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd0,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b4e_blk00000b4f_sig0000145f,
      Q31 => NLW_blk00000001_blk00000b4e_blk00000b4f_blk00000b52_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b4e_blk00000b4f_sig0000145e,
      A(3) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(2) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(1) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d,
      A(0) => blk00000001_blk00000b4e_blk00000b4f_sig0000145d
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b51 : VCC
    port map (
      P => blk00000001_blk00000b4e_blk00000b4f_sig0000145e
    );
  blk00000001_blk00000b4e_blk00000b4f_blk00000b50 : GND
    port map (
      G => blk00000001_blk00000b4e_blk00000b4f_sig0000145d
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b65 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b5a_blk00000b5b_sig0000147d,
      Q => blk00000001_sig00000db2
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b64 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd6,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b5a_blk00000b5b_sig0000147d,
      Q31 => NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b64_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b5a_blk00000b5b_sig00001479,
      A(3) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(2) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(1) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(0) => blk00000001_blk00000b5a_blk00000b5b_sig00001478
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b63 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b5a_blk00000b5b_sig0000147c,
      Q => blk00000001_sig00000db1
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b62 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd5,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b5a_blk00000b5b_sig0000147c,
      Q31 => NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b62_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b5a_blk00000b5b_sig00001479,
      A(3) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(2) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(1) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(0) => blk00000001_blk00000b5a_blk00000b5b_sig00001478
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b61 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b5a_blk00000b5b_sig0000147b,
      Q => blk00000001_sig00000db0
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b60 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd4,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b5a_blk00000b5b_sig0000147b,
      Q31 => NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b60_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b5a_blk00000b5b_sig00001479,
      A(3) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(2) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(1) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(0) => blk00000001_blk00000b5a_blk00000b5b_sig00001478
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b5f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b5a_blk00000b5b_sig0000147a,
      Q => blk00000001_sig00000daf
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b5e : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd9,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b5a_blk00000b5b_sig0000147a,
      Q31 => NLW_blk00000001_blk00000b5a_blk00000b5b_blk00000b5e_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b5a_blk00000b5b_sig00001479,
      A(3) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(2) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(1) => blk00000001_blk00000b5a_blk00000b5b_sig00001478,
      A(0) => blk00000001_blk00000b5a_blk00000b5b_sig00001478
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b5d : VCC
    port map (
      P => blk00000001_blk00000b5a_blk00000b5b_sig00001479
    );
  blk00000001_blk00000b5a_blk00000b5b_blk00000b5c : GND
    port map (
      G => blk00000001_blk00000b5a_blk00000b5b_sig00001478
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b71 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b66_blk00000b67_sig00001498,
      Q => blk00000001_sig00000dae
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b70 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd8,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b66_blk00000b67_sig00001498,
      Q31 => NLW_blk00000001_blk00000b66_blk00000b67_blk00000b70_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b66_blk00000b67_sig00001494,
      A(3) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(2) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(1) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(0) => blk00000001_blk00000b66_blk00000b67_sig00001493
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b66_blk00000b67_sig00001497,
      Q => blk00000001_sig00000dad
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6e : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd2,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b66_blk00000b67_sig00001497,
      Q31 => NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6e_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b66_blk00000b67_sig00001494,
      A(3) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(2) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(1) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(0) => blk00000001_blk00000b66_blk00000b67_sig00001493
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b66_blk00000b67_sig00001496,
      Q => blk00000001_sig00000dac
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6c : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd7,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b66_blk00000b67_sig00001496,
      Q31 => NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6c_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b66_blk00000b67_sig00001494,
      A(3) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(2) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(1) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(0) => blk00000001_blk00000b66_blk00000b67_sig00001493
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b66_blk00000b67_sig00001495,
      Q => blk00000001_sig00000dab
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b6a : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd0,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b66_blk00000b67_sig00001495,
      Q31 => NLW_blk00000001_blk00000b66_blk00000b67_blk00000b6a_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b66_blk00000b67_sig00001494,
      A(3) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(2) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(1) => blk00000001_blk00000b66_blk00000b67_sig00001493,
      A(0) => blk00000001_blk00000b66_blk00000b67_sig00001493
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b69 : VCC
    port map (
      P => blk00000001_blk00000b66_blk00000b67_sig00001494
    );
  blk00000001_blk00000b66_blk00000b67_blk00000b68 : GND
    port map (
      G => blk00000001_blk00000b66_blk00000b67_sig00001493
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b7d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b72_blk00000b73_sig000014b3,
      Q => blk00000001_sig00000daa
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b7c : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000ddb,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b72_blk00000b73_sig000014b3,
      Q31 => NLW_blk00000001_blk00000b72_blk00000b73_blk00000b7c_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b72_blk00000b73_sig000014af,
      A(3) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(2) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(1) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(0) => blk00000001_blk00000b72_blk00000b73_sig000014ae
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b7b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b72_blk00000b73_sig000014b2,
      Q => blk00000001_sig00000da9
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b7a : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd5,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b72_blk00000b73_sig000014b2,
      Q31 => NLW_blk00000001_blk00000b72_blk00000b73_blk00000b7a_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b72_blk00000b73_sig000014af,
      A(3) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(2) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(1) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(0) => blk00000001_blk00000b72_blk00000b73_sig000014ae
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b79 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b72_blk00000b73_sig000014b1,
      Q => blk00000001_sig00000da8
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b78 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dda,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b72_blk00000b73_sig000014b1,
      Q31 => NLW_blk00000001_blk00000b72_blk00000b73_blk00000b78_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b72_blk00000b73_sig000014af,
      A(3) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(2) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(1) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(0) => blk00000001_blk00000b72_blk00000b73_sig000014ae
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b77 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000008e,
      D => blk00000001_blk00000b72_blk00000b73_sig000014b0,
      Q => blk00000001_sig00000da7
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b76 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_sig00000dd9,
      CE => blk00000001_sig0000008e,
      Q => blk00000001_blk00000b72_blk00000b73_sig000014b0,
      Q31 => NLW_blk00000001_blk00000b72_blk00000b73_blk00000b76_Q31_UNCONNECTED,
      A(4) => blk00000001_blk00000b72_blk00000b73_sig000014af,
      A(3) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(2) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(1) => blk00000001_blk00000b72_blk00000b73_sig000014ae,
      A(0) => blk00000001_blk00000b72_blk00000b73_sig000014ae
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b75 : VCC
    port map (
      P => blk00000001_blk00000b72_blk00000b73_sig000014af
    );
  blk00000001_blk00000b72_blk00000b73_blk00000b74 : GND
    port map (
      G => blk00000001_blk00000b72_blk00000b73_sig000014ae
    );

end STRUCTURE;

-- synthesis translate_on

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity axi_sgiface is
    generic (
        -- AXI specific.
        -- TODO: need to figure out a way to pass these generics from outside
        C_S_AXI_SUPPORT_BURST   : integer := 0;
        -- TODO: fix the internal ID width to 8
        C_S_AXI_ID_WIDTH        : integer := 8;
        C_S_AXI_DATA_WIDTH      : integer := 32;
        C_S_AXI_ADDR_WIDTH      : integer := 32;
        C_S_AXI_TOTAL_ADDR_LEN  : integer := 12;
        C_S_AXI_LINEAR_ADDR_LEN : integer := 8;
        C_S_AXI_BANK_ADDR_LEN   : integer := 2;
        C_S_AXI_AWLEN_WIDTH     : integer := 8;
        C_S_AXI_ARLEN_WIDTH     : integer := 8
    );
    port (
        -- General.
        AXI_AClk      : in  std_logic;
        AXI_AResetN    : in  std_logic;
        -- not used
        AXI_Ce        : in  std_logic;
  
        -- AXI Port.
        S_AXI_AWADDR  : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_AWID    : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_AWLEN   : in  std_logic_vector(C_S_AXI_AWLEN_WIDTH-1 downto 0);
        S_AXI_AWSIZE  : in  std_logic_vector(2 downto 0);
        S_AXI_AWBURST : in  std_logic_vector(1 downto 0);
        S_AXI_AWLOCK  : in  std_logic_vector(1 downto 0);
        S_AXI_AWCACHE : in  std_logic_vector(3 downto 0);
        S_AXI_AWPROT  : in  std_logic_vector(2 downto 0);
        S_AXI_AWVALID : in  std_logic;
        S_AXI_AWREADY : out std_logic;
        
        S_AXI_WLAST   : in  std_logic;
        S_AXI_WDATA   : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_WSTRB   : in  std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
        S_AXI_WVALID  : in  std_logic;
        S_AXI_WREADY  : out std_logic;
        
        S_AXI_BRESP   : out std_logic_vector(1 downto 0);
        S_AXI_BID     : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_BVALID  : out std_logic;
        S_AXI_BREADY  : in  std_logic;
        
        S_AXI_ARADDR  : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_ARID    : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_ARLEN   : in  std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
        S_AXI_ARSIZE  : in  std_logic_vector(2 downto 0);
        S_AXI_ARBURST : in  std_logic_vector(1 downto 0);
        S_AXI_ARLOCK  : in  std_logic_vector(1 downto 0);
        S_AXI_ARCACHE : in  std_logic_vector(3 downto 0);
        S_AXI_ARPROT  : in  std_logic_vector(2 downto 0);
        S_AXI_ARVALID : in  std_logic;
        S_AXI_ARREADY : out std_logic;
        
        -- 'From Register'
        -- 'STATUS'
        sm_STATUS_dout : in std_logic_vector(32-1 downto 0);
        -- 'To Register'
        -- 'Timing'
        sm_Timing_dout : in std_logic_vector(32-1 downto 0);
        sm_Timing_din  : out std_logic_vector(32-1 downto 0);
        sm_Timing_en   : out std_logic;
        -- 'Config'
        sm_Config_dout : in std_logic_vector(32-1 downto 0);
        sm_Config_din  : out std_logic_vector(32-1 downto 0);
        sm_Config_en   : out std_logic;
        -- 'PKT_BUF_SEL'
        sm_PKT_BUF_SEL_dout : in std_logic_vector(32-1 downto 0);
        sm_PKT_BUF_SEL_din  : out std_logic_vector(32-1 downto 0);
        sm_PKT_BUF_SEL_en   : out std_logic;
        -- 'Output_Scaling'
        sm_Output_Scaling_dout : in std_logic_vector(32-1 downto 0);
        sm_Output_Scaling_din  : out std_logic_vector(32-1 downto 0);
        sm_Output_Scaling_en   : out std_logic;
        -- 'TX_START'
        sm_TX_START_dout : in std_logic_vector(32-1 downto 0);
        sm_TX_START_din  : out std_logic_vector(32-1 downto 0);
        sm_TX_START_en   : out std_logic;
        -- 'FFT_Config'
        sm_FFT_Config_dout : in std_logic_vector(32-1 downto 0);
        sm_FFT_Config_din  : out std_logic_vector(32-1 downto 0);
        sm_FFT_Config_en   : out std_logic;
        -- 'From FIFO'
        -- 'To FIFO'
        -- 'Shared Memory'

        S_AXI_RLAST   : out std_logic;
        S_AXI_RID     : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_RDATA   : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_RRESP   : out std_logic_vector(1 downto 0);
        S_AXI_RVALID  : out std_logic;
        S_AXI_RREADY  : in  std_logic
    );
end entity axi_sgiface;

architecture IMP of axi_sgiface is

-- Internal signals for write channel.
signal S_AXI_BVALID_i       : std_logic;
signal S_AXI_BID_i          : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
signal S_AXI_WREADY_i       : std_logic;
  
-- Internal signals for read channels.
signal S_AXI_ARLEN_i        : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
signal S_AXI_RLAST_i        : std_logic;
signal S_AXI_RREADY_i       : std_logic;
signal S_AXI_RVALID_i       : std_logic;
signal S_AXI_RDATA_i        : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal S_AXI_RID_i          : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);

-- for read channel
signal read_bank_addr_i     : std_logic_vector(C_S_AXI_BANK_ADDR_LEN-1 downto 0);
signal read_linear_addr_i   : std_logic_vector(C_S_AXI_LINEAR_ADDR_LEN-1 downto 0);
-- for write channel
signal write_bank_addr_i    : std_logic_vector(C_S_AXI_BANK_ADDR_LEN-1 downto 0);
signal write_linear_addr_i  : std_logic_vector(C_S_AXI_LINEAR_ADDR_LEN-1 downto 0);

signal reg_bank_out_i       : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal fifo_bank_out_i      : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal shmem_bank_out_i     : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    
-- 'From Register'
-- 'STATUS'
signal sm_STATUS_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'To Register'
-- 'Timing'
signal sm_Timing_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Timing_en_i    : std_logic;
signal sm_Timing_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'Config'
signal sm_Config_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Config_en_i    : std_logic;
signal sm_Config_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'PKT_BUF_SEL'
signal sm_PKT_BUF_SEL_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_PKT_BUF_SEL_en_i    : std_logic;
signal sm_PKT_BUF_SEL_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'Output_Scaling'
signal sm_Output_Scaling_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Output_Scaling_en_i    : std_logic;
signal sm_Output_Scaling_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'TX_START'
signal sm_TX_START_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_TX_START_en_i    : std_logic;
signal sm_TX_START_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'FFT_Config'
signal sm_FFT_Config_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_FFT_Config_en_i    : std_logic;
signal sm_FFT_Config_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'From FIFO'
-- 'To FIFO'
-- 'Shared Memory'

type t_read_state is (IDLE, READ_PREP, READ_DATA);
signal read_state : t_read_state;

type t_write_state is (IDLE, WRITE_DATA, WRITE_RESPONSE);
signal write_state : t_write_state;

type t_memmap_state is (READ, WRITE);
signal memmap_state : t_memmap_state;

constant C_READ_PREP_DELAY : std_logic_vector(1 downto 0) := "11";

signal read_prep_counter : std_logic_vector(1 downto 0);
signal read_addr_counter : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
signal read_data_counter : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);

-- enable of shared BRAMs
signal s_shram_en : std_logic;

signal write_addr_valid : std_logic;
signal write_ready : std_logic;

-- 're' of From/To FIFOs
signal s_fifo_re : std_logic;
-- 'we' of To FIFOs
signal s_fifo_we : std_logic;

begin

-- enable for 'Shared Memory' blocks

-- conversion to match with the data bus width
-- 'From Register'
-- 'STATUS'
gen_sm_STATUS_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_STATUS_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_STATUS_dout_i;
sm_STATUS_dout_i(32-1 downto 0) <= sm_STATUS_dout;
-- 'To Register'
-- 'Timing'
sm_Timing_din     <= sm_Timing_din_i(32-1 downto 0);
sm_Timing_en      <= sm_Timing_en_i;
gen_sm_Timing_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Timing_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Timing_dout_i;
sm_Timing_dout_i(32-1 downto 0) <= sm_Timing_dout;
-- 'Config'
sm_Config_din     <= sm_Config_din_i(32-1 downto 0);
sm_Config_en      <= sm_Config_en_i;
gen_sm_Config_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Config_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Config_dout_i;
sm_Config_dout_i(32-1 downto 0) <= sm_Config_dout;
-- 'PKT_BUF_SEL'
sm_PKT_BUF_SEL_din     <= sm_PKT_BUF_SEL_din_i(32-1 downto 0);
sm_PKT_BUF_SEL_en      <= sm_PKT_BUF_SEL_en_i;
gen_sm_PKT_BUF_SEL_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_PKT_BUF_SEL_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_PKT_BUF_SEL_dout_i;
sm_PKT_BUF_SEL_dout_i(32-1 downto 0) <= sm_PKT_BUF_SEL_dout;
-- 'Output_Scaling'
sm_Output_Scaling_din     <= sm_Output_Scaling_din_i(32-1 downto 0);
sm_Output_Scaling_en      <= sm_Output_Scaling_en_i;
gen_sm_Output_Scaling_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Output_Scaling_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Output_Scaling_dout_i;
sm_Output_Scaling_dout_i(32-1 downto 0) <= sm_Output_Scaling_dout;
-- 'TX_START'
sm_TX_START_din     <= sm_TX_START_din_i(32-1 downto 0);
sm_TX_START_en      <= sm_TX_START_en_i;
gen_sm_TX_START_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_TX_START_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_TX_START_dout_i;
sm_TX_START_dout_i(32-1 downto 0) <= sm_TX_START_dout;
-- 'FFT_Config'
sm_FFT_Config_din     <= sm_FFT_Config_din_i(32-1 downto 0);
sm_FFT_Config_en      <= sm_FFT_Config_en_i;
gen_sm_FFT_Config_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_FFT_Config_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_FFT_Config_dout_i;
sm_FFT_Config_dout_i(32-1 downto 0) <= sm_FFT_Config_dout;
-- 'From FIFO'
-- 'To FIFO'
-- 'Shared Memory'

ReadWriteSelect: process(memmap_state) is begin
    if (memmap_state = READ) then
    else
    end if;
end process ReadWriteSelect;

-----------------------------------------------------------------------------
-- address for 'Shared Memory'
-----------------------------------------------------------------------------
SharedMemory_Addr_ResetN : process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            memmap_state <= READ;
        else
            if (S_AXI_AWVALID = '1') then
                -- write operation
                memmap_state <= WRITE;
            elsif (S_AXI_ARVALID = '1') then
                -- read operation
                memmap_state <= READ;
            end if;
        end if;
    end if;
end process SharedMemory_Addr_ResetN;

-----------------------------------------------------------------------------
-- WRITE Command Control
-----------------------------------------------------------------------------
S_AXI_BID     <= S_AXI_BID_i;
S_AXI_BVALID  <= S_AXI_BVALID_i;
S_AXI_WREADY  <= S_AXI_WREADY_i;
-- No error checking
S_AXI_BRESP  <= (others=>'0');

PROC_AWREADY_ACK: process(read_state, write_state, S_AXI_ARVALID, S_AXI_AWVALID) is begin
    if (write_state = IDLE and S_AXI_AWVALID = '1' and read_state = IDLE) then
        S_AXI_AWREADY <= S_AXI_AWVALID;
    else
        S_AXI_AWREADY <= '0';
    end if;
end process PROC_AWREADY_ACK;

Cmd_Decode_Write: process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            write_addr_valid    <= '0';
            write_ready         <= '0';
            s_fifo_we           <= '0';
            S_AXI_BVALID_i      <= '0';
            S_AXI_BID_i         <= (others => '0');
            write_bank_addr_i   <= (others => '0');
            write_linear_addr_i <= (others => '0');
        else
            if (write_state = IDLE) then
                if (S_AXI_AWVALID = '1' and read_state = IDLE) then
                    -- reflect awid
                    S_AXI_BID_i <= S_AXI_AWID;

                    -- latch bank and linear addresses
                    write_bank_addr_i   <= S_AXI_AWADDR(C_S_AXI_TOTAL_ADDR_LEN-1 downto C_S_AXI_LINEAR_ADDR_LEN+2);
                    write_linear_addr_i <= S_AXI_AWADDR(C_S_AXI_LINEAR_ADDR_LEN+1 downto 2);
                    write_addr_valid <= '1';
                    s_fifo_we <= '1';

                    -- write state transition
                    write_state <= WRITE_DATA;
                end if;
            elsif (write_state = WRITE_DATA) then
                write_ready <= '1';
                s_fifo_we <= '0';
                write_addr_valid <= S_AXI_WVALID;
                
                if (S_AXI_WVALID = '1' and write_ready = '1') then
                    write_linear_addr_i <= Std_Logic_Vector(unsigned(write_linear_addr_i) + 1);
                end if;

                if (S_AXI_WLAST = '1' and write_ready = '1') then
                    -- start responding through B channel upon the last write data sample
                    S_AXI_BVALID_i <= '1';
                    -- write data is over
                    write_addr_valid <= '0';
                    write_ready <= '0';
                    -- write state transition
                    write_state <= WRITE_RESPONSE;
                end if;
            elsif (write_state = WRITE_RESPONSE) then

                if (S_AXI_BREADY = '1') then
                    -- write respond is over
                    S_AXI_BVALID_i <= '0';
                    S_AXI_BID_i <= (others => '0');

                    -- write state transition
                    write_state <= IDLE;
                end if;
            end if;
        end if;
    end if;
end process Cmd_Decode_Write;

Write_Linear_Addr_Decode : process(AXI_AClk) is 

begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            -- 'To Register'
            -- Timing din/en
            sm_Timing_din_i <= (others => '0');
            sm_Timing_en_i <= '0';
            -- Config din/en
            sm_Config_din_i <= (others => '0');
            sm_Config_en_i <= '0';
            -- PKT_BUF_SEL din/en
            sm_PKT_BUF_SEL_din_i <= (others => '0');
            sm_PKT_BUF_SEL_en_i <= '0';
            -- Output_Scaling din/en
            sm_Output_Scaling_din_i <= (others => '0');
            sm_Output_Scaling_en_i <= '0';
            -- TX_START din/en
            sm_TX_START_din_i <= (others => '0');
            sm_TX_START_en_i <= '0';
            -- FFT_Config din/en
            sm_FFT_Config_din_i <= (others => '0');
            sm_FFT_Config_en_i <= '0';
            -- 'To FIFO'
            -- 'Shared Memory'
        else
            -- default assignments

            -- 'To Register'
            if (unsigned(write_bank_addr_i) = 2) then
                if (unsigned(write_linear_addr_i) = 0) then
                    -- Timing din/en
                    sm_Timing_din_i <= S_AXI_WDATA;
                    sm_Timing_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 1) then
                    -- Config din/en
                    sm_Config_din_i <= S_AXI_WDATA;
                    sm_Config_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 2) then
                    -- PKT_BUF_SEL din/en
                    sm_PKT_BUF_SEL_din_i <= S_AXI_WDATA;
                    sm_PKT_BUF_SEL_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 3) then
                    -- Output_Scaling din/en
                    sm_Output_Scaling_din_i <= S_AXI_WDATA;
                    sm_Output_Scaling_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 4) then
                    -- TX_START din/en
                    sm_TX_START_din_i <= S_AXI_WDATA;
                    sm_TX_START_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 5) then
                    -- FFT_Config din/en
                    sm_FFT_Config_din_i <= S_AXI_WDATA;
                    sm_FFT_Config_en_i  <= write_addr_valid;
                end if;
            end if;        
        
        
        end if;
    end if;
end process Write_Linear_Addr_Decode;
 
-----------------------------------------------------------------------------
-- READ Control
-----------------------------------------------------------------------------

S_AXI_RDATA  <= S_AXI_RDATA_i;
S_AXI_RVALID  <= S_AXI_RVALID_i;
S_AXI_RLAST   <= S_AXI_RLAST_i;
S_AXI_RID     <= S_AXI_RID_i;
-- TODO: no error checking
S_AXI_RRESP <= (others=>'0');

PROC_ARREADY_ACK: process(read_state, S_AXI_ARVALID, write_state, S_AXI_AWVALID) is begin
    -- Note: WRITE has higher priority than READ
    if (read_state = IDLE and S_AXI_ARVALID = '1' and write_state = IDLE and S_AXI_AWVALID /= '1') then
        S_AXI_ARREADY <= S_AXI_ARVALID;
    else
        S_AXI_ARREADY <= '0';
    end if;
end process PROC_ARREADY_ACK;

S_AXI_WREADY_i <= write_ready;

Process_Sideband: process(write_state, read_state) is begin
    if (read_state = READ_PREP) then
        s_shram_en <= '1';
    elsif (read_state = READ_DATA) then
        s_shram_en <= S_AXI_RREADY;
    elsif (write_state = WRITE_DATA) then
        s_shram_en <= S_AXI_WVALID;
    else
        s_shram_en <= '0';
    end if;
end process Process_Sideband;

Cmd_Decode_Read: process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            S_AXI_RVALID_i <= '0';
            read_bank_addr_i    <= (others => '0');
            read_linear_addr_i  <= (others => '0');
            S_AXI_ARLEN_i       <= (others => '0');
            S_AXI_RLAST_i       <= '0';
            S_AXI_RID_i         <= (others => '0');
            read_state          <= IDLE;
            read_prep_counter   <= (others => '0');
            read_addr_counter   <= (others => '0');
            read_data_counter   <= (others => '0');
        else
            -- default assignments
            s_fifo_re <= '0';

            if (read_state = IDLE) then
                -- Note WRITE has higher priority than READ
                if (S_AXI_ARVALID = '1' and write_state = IDLE and S_AXI_AWVALID /= '1') then
                    -- extract bank and linear addresses
                    read_bank_addr_i    <= S_AXI_ARADDR(C_S_AXI_TOTAL_ADDR_LEN-1 downto C_S_AXI_LINEAR_ADDR_LEN+2);
                    read_linear_addr_i  <= S_AXI_ARADDR(C_S_AXI_LINEAR_ADDR_LEN+1 downto 2);
                    s_fifo_re <= '1';

                    -- reflect arid
                    S_AXI_RID_i <= S_AXI_ARID;

                    -- load read liner address and data counter
                    read_addr_counter <= S_AXI_ARLEN;
                    read_data_counter <= S_AXI_ARLEN;

                    -- load read preparation counter
                    read_prep_counter <= C_READ_PREP_DELAY;
                    -- read state transition
                    read_state <= READ_PREP;
                end if;
            elsif (read_state = READ_PREP) then
                if (unsigned(read_prep_counter) = 0) then
                    if (unsigned(read_data_counter) = 0) then
                        -- tag the last data generated by the slave
                        S_AXI_RLAST_i <= '1';
                    end if;
                    -- valid data appears
                    S_AXI_RVALID_i <= '1';
                    -- read state transition
                    read_state <= READ_DATA;
                else
                    -- decrease read preparation counter
                    read_prep_counter <= Std_Logic_Vector(unsigned(read_prep_counter) - 1);
                end if;

                if (unsigned(read_prep_counter) /= 3 and unsigned(read_addr_counter) /= 0) then
                    -- decrease address counter
                    read_addr_counter <= Std_Logic_Vector(unsigned(read_addr_counter) - 1);
                    -- increase linear address (no band crossing)
                    read_linear_addr_i <= Std_Logic_Vector(unsigned(read_linear_addr_i) + 1);
                end if;
            elsif (read_state = READ_DATA) then
                if (S_AXI_RREADY = '1') then
                    if (unsigned(read_data_counter) = 1) then
                        -- tag the last data generated by the slave
                        S_AXI_RLAST_i <= '1';
                    end if;

                    if (unsigned(read_data_counter) = 0) then
                        -- arid
                        S_AXI_RID_i <= (others => '0');
                        -- rlast
                        S_AXI_RLAST_i <= '0';
                        -- no more valid data
                        S_AXI_RVALID_i <= '0';
                        -- read state transition
                        read_state <= IDLE;
                    else
                        -- decrease read preparation counter
                        read_data_counter <= Std_Logic_Vector(unsigned(read_data_counter) - 1);

                        if (unsigned(read_addr_counter) /= 0) then
                            -- decrease address counter
                            read_addr_counter <= Std_Logic_Vector(unsigned(read_addr_counter) - 1);
                            -- increase linear address (no band crossing)
                            read_linear_addr_i <= Std_Logic_Vector(unsigned(read_linear_addr_i) + 1);
                        end if;
                    end if;
                end if;
            end if;

        end if;
    end if;
end process Cmd_Decode_Read;

Read_Linear_Addr_Decode : process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            reg_bank_out_i   <= (others => '0');
            fifo_bank_out_i  <= (others => '0');
            shmem_bank_out_i <= (others => '0');
            S_AXI_RDATA_i    <= (others => '0');
        else
            if (unsigned(read_bank_addr_i) = 2) then
                -- 'From Register'
                if (unsigned(read_linear_addr_i) = 6) then
                    -- 'STATUS' dout
                    reg_bank_out_i <= sm_STATUS_dout_i;
                end if;
                -- 'To Register' (with register readback)
                if (unsigned(read_linear_addr_i) = 0) then
                    -- 'Timing' dout
                    reg_bank_out_i <= sm_Timing_dout_i;
                elsif (unsigned(read_linear_addr_i) = 1) then
                    -- 'Config' dout
                    reg_bank_out_i <= sm_Config_dout_i;
                elsif (unsigned(read_linear_addr_i) = 2) then
                    -- 'PKT_BUF_SEL' dout
                    reg_bank_out_i <= sm_PKT_BUF_SEL_dout_i;
                elsif (unsigned(read_linear_addr_i) = 3) then
                    -- 'Output_Scaling' dout
                    reg_bank_out_i <= sm_Output_Scaling_dout_i;
                elsif (unsigned(read_linear_addr_i) = 4) then
                    -- 'TX_START' dout
                    reg_bank_out_i <= sm_TX_START_dout_i;
                elsif (unsigned(read_linear_addr_i) = 5) then
                    -- 'FFT_Config' dout
                    reg_bank_out_i <= sm_FFT_Config_dout_i;
                end if;

                S_AXI_RDATA_i <= reg_bank_out_i;
            elsif (unsigned(read_bank_addr_i) = 1) then
                -- 'From FIFO'
                -- 'To FIFO'

                S_AXI_RDATA_i <= fifo_bank_out_i;
            elsif (unsigned(read_bank_addr_i) = 0 and s_shram_en = '1') then
                -- 'Shared Memory'

                S_AXI_RDATA_i <= shmem_bank_out_i;
            end if;
        end if;
    end if;
end process Read_Linear_Addr_Decode;

end architecture IMP;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_0d20f96564 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_0d20f96564;


architecture behavior of concat_0d20f96564 is
  signal in0_1_23: boolean;
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= ((in0) = "1");
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(boolean_to_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c462ec0feb is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c462ec0feb;


architecture behavior of constant_c462ec0feb is
begin
  op <= "111111";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlcounter_free_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free_wlan_phy_tx_pmd ;
architecture behavior of xlcounter_free_wlan_phy_tx_pmd is
  component cntr_11_0_f068fb73312ae1e5
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_f068fb73312ae1e5:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_f068fb73312ae1e5:
    component is "true";
  attribute box_type of cntr_11_0_f068fb73312ae1e5:
    component  is "black_box";
  component cntr_11_0_86806e294f737f4c
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_86806e294f737f4c:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_86806e294f737f4c:
    component is "true";
  attribute box_type of cntr_11_0_86806e294f737f4c:
    component  is "black_box";
  component cntr_11_0_511eb7a1af6f3f2a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_511eb7a1af6f3f2a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_511eb7a1af6f3f2a:
    component is "true";
  attribute box_type of cntr_11_0_511eb7a1af6f3f2a:
    component  is "black_box";
  component cntr_11_0_d5912692bc2e79ac
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d5912692bc2e79ac:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d5912692bc2e79ac:
    component is "true";
  attribute box_type of cntr_11_0_d5912692bc2e79ac:
    component  is "black_box";
  component cntr_11_0_36e2bb554c95560d
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_36e2bb554c95560d:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_36e2bb554c95560d:
    component is "true";
  attribute box_type of cntr_11_0_36e2bb554c95560d:
    component  is "black_box";
  component cntr_11_0_87d991c7bcfe987f
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_87d991c7bcfe987f:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_87d991c7bcfe987f:
    component is "true";
  attribute box_type of cntr_11_0_87d991c7bcfe987f:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_f068fb73312ae1e5")) generate
    core_instance0: cntr_11_0_f068fb73312ae1e5
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_86806e294f737f4c")) generate
    core_instance1: cntr_11_0_86806e294f737f4c
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp2: if ((core_name0 = "cntr_11_0_511eb7a1af6f3f2a")) generate
    core_instance2: cntr_11_0_511eb7a1af6f3f2a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp3: if ((core_name0 = "cntr_11_0_d5912692bc2e79ac")) generate
    core_instance3: cntr_11_0_d5912692bc2e79ac
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp4: if ((core_name0 = "cntr_11_0_36e2bb554c95560d")) generate
    core_instance4: cntr_11_0_36e2bb554c95560d
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp5: if ((core_name0 = "cntr_11_0_87d991c7bcfe987f")) generate
    core_instance5: cntr_11_0_87d991c7bcfe987f
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer :=  0;
           reset        : integer :=  0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        rst     : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if ((reg_retiming = 0) and (reset = 0)) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if ((reg_retiming = 1) or (reset = 1)) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => rst,
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_dist_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    addr_width: integer := 2;
    latency: integer := 0;
    c_width: integer := 12;
    c_address_width: integer := 4
  );
  port (
    addr: in std_logic_vector(addr_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_dist_wlan_phy_tx_pmd ;
architecture behavior of xlsprom_dist_wlan_phy_tx_pmd is
  component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i           : in std_logic_vector(width - 1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width - 1 downto 0));
  end component;
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  constant num_extra_addr_bits: integer := (c_address_width - addr_width);
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_ce: std_logic;
  component dmg_72_48a0132db6517610
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_48a0132db6517610:
    component is true;
  attribute fpga_dont_touch of dmg_72_48a0132db6517610:
    component is "true";
  attribute box_type of dmg_72_48a0132db6517610:
    component  is "black_box";
  component dmg_72_2be916f69ff4e5b8
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_2be916f69ff4e5b8:
    component is true;
  attribute fpga_dont_touch of dmg_72_2be916f69ff4e5b8:
    component is "true";
  attribute box_type of dmg_72_2be916f69ff4e5b8:
    component  is "black_box";
  component dmg_72_58f1077b49388e77
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_58f1077b49388e77:
    component is true;
  attribute fpga_dont_touch of dmg_72_58f1077b49388e77:
    component is "true";
  attribute box_type of dmg_72_58f1077b49388e77:
    component  is "black_box";
  component dmg_72_d59da422e431313e
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_d59da422e431313e:
    component is true;
  attribute fpga_dont_touch of dmg_72_d59da422e431313e:
    component is "true";
  attribute box_type of dmg_72_d59da422e431313e:
    component  is "black_box";
  component dmg_72_134e91999cae8947
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_134e91999cae8947:
    component is true;
  attribute fpga_dont_touch of dmg_72_134e91999cae8947:
    component is "true";
  attribute box_type of dmg_72_134e91999cae8947:
    component  is "black_box";
  component dmg_72_06262d82a068201e
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_06262d82a068201e:
    component is true;
  attribute fpga_dont_touch of dmg_72_06262d82a068201e:
    component is "true";
  attribute box_type of dmg_72_06262d82a068201e:
    component  is "black_box";
  component dmg_72_d16d082a6bc00ceb
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_d16d082a6bc00ceb:
    component is true;
  attribute fpga_dont_touch of dmg_72_d16d082a6bc00ceb:
    component is "true";
  attribute box_type of dmg_72_d16d082a6bc00ceb:
    component  is "black_box";
  component dmg_72_2b0650236539a42c
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_2b0650236539a42c:
    component is true;
  attribute fpga_dont_touch of dmg_72_2b0650236539a42c:
    component is "true";
  attribute box_type of dmg_72_2b0650236539a42c:
    component  is "black_box";
begin
  need_to_pad_addr: if num_extra_addr_bits > 0 generate
      core_addr(c_address_width - 1 downto addr_width) <= (others => '0');
    core_addr(addr_width - 1 downto 0) <= addr;
  end generate;
  no_need_to_pad_addr: if num_extra_addr_bits = 0 generate
    core_addr <= addr;
  end generate;
  core_ce <= ce and en(0);
  comp0: if ((core_name0 = "dmg_72_48a0132db6517610")) generate
    core_instance0: dmg_72_48a0132db6517610
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  comp1: if ((core_name0 = "dmg_72_2be916f69ff4e5b8")) generate
    core_instance1: dmg_72_2be916f69ff4e5b8
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  comp2: if ((core_name0 = "dmg_72_58f1077b49388e77")) generate
    core_instance2: dmg_72_58f1077b49388e77
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp3: if ((core_name0 = "dmg_72_d59da422e431313e")) generate
    core_instance3: dmg_72_d59da422e431313e
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp4: if ((core_name0 = "dmg_72_134e91999cae8947")) generate
    core_instance4: dmg_72_134e91999cae8947
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp5: if ((core_name0 = "dmg_72_06262d82a068201e")) generate
    core_instance5: dmg_72_06262d82a068201e
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp6: if ((core_name0 = "dmg_72_d16d082a6bc00ceb")) generate
    core_instance6: dmg_72_d16d082a6bc00ceb
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  comp7: if ((core_name0 = "dmg_72_2b0650236539a42c")) generate
    core_instance7: dmg_72_2b0650236539a42c
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_0_or_1: if (latency <= 1)
  generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_80f90b97d0 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_80f90b97d0;


architecture behavior of logical_80f90b97d0 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mcode_block_00412594a7 is
  port (
    sym_cfg : in std_logic_vector((18 - 1) downto 0);
    load_base_rate : out std_logic_vector((1 - 1) downto 0);
    rotate_bpsk : out std_logic_vector((1 - 1) downto 0);
    load_htstf : out std_logic_vector((1 - 1) downto 0);
    load_htltf : out std_logic_vector((1 - 1) downto 0);
    load_full_rate : out std_logic_vector((1 - 1) downto 0);
    pilot_shift : out std_logic_vector((2 - 1) downto 0);
    cyclic_prefix : out std_logic_vector((5 - 1) downto 0);
    cyclic_shift : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mcode_block_00412594a7;


architecture behavior of mcode_block_00412594a7 is
  signal sym_cfg_1_142: unsigned((18 - 1) downto 0);
  signal slice_19_26: unsigned((1 - 1) downto 0);
  signal load_base_rate_19_1_rel: boolean;
  signal slice_20_26: unsigned((1 - 1) downto 0);
  signal rotate_bpsk_20_1_rel: boolean;
  signal slice_21_26: unsigned((1 - 1) downto 0);
  signal load_htstf_21_1_rel: boolean;
  signal slice_22_26: unsigned((1 - 1) downto 0);
  signal load_htltf_22_1_rel: boolean;
  signal slice_23_26: unsigned((1 - 1) downto 0);
  signal load_full_rate_23_1_rel: boolean;
  signal pilot_shift_24_1_slice: unsigned((2 - 1) downto 0);
  signal cyclic_prefix_26_1_slice: unsigned((5 - 1) downto 0);
  signal cyclic_shift_27_1_slice: unsigned((3 - 1) downto 0);
begin
  sym_cfg_1_142 <= std_logic_vector_to_unsigned(sym_cfg);
  slice_19_26 <= u2u_slice(sym_cfg_1_142, 0, 0);
  load_base_rate_19_1_rel <= slice_19_26 = std_logic_vector_to_unsigned("1");
  slice_20_26 <= u2u_slice(sym_cfg_1_142, 1, 1);
  rotate_bpsk_20_1_rel <= slice_20_26 = std_logic_vector_to_unsigned("1");
  slice_21_26 <= u2u_slice(sym_cfg_1_142, 2, 2);
  load_htstf_21_1_rel <= slice_21_26 = std_logic_vector_to_unsigned("1");
  slice_22_26 <= u2u_slice(sym_cfg_1_142, 3, 3);
  load_htltf_22_1_rel <= slice_22_26 = std_logic_vector_to_unsigned("1");
  slice_23_26 <= u2u_slice(sym_cfg_1_142, 4, 4);
  load_full_rate_23_1_rel <= slice_23_26 = std_logic_vector_to_unsigned("1");
  pilot_shift_24_1_slice <= u2u_slice(sym_cfg_1_142, 6, 5);
  cyclic_prefix_26_1_slice <= u2u_slice(sym_cfg_1_142, 12, 8);
  cyclic_shift_27_1_slice <= u2u_slice(sym_cfg_1_142, 15, 13);
  load_base_rate <= boolean_to_vector(load_base_rate_19_1_rel);
  rotate_bpsk <= boolean_to_vector(rotate_bpsk_20_1_rel);
  load_htstf <= boolean_to_vector(load_htstf_21_1_rel);
  load_htltf <= boolean_to_vector(load_htltf_22_1_rel);
  load_full_rate <= boolean_to_vector(load_full_rate_23_1_rel);
  pilot_shift <= unsigned_to_std_logic_vector(pilot_shift_24_1_slice);
  cyclic_prefix <= unsigned_to_std_logic_vector(cyclic_prefix_26_1_slice);
  cyclic_shift <= unsigned_to_std_logic_vector(cyclic_shift_27_1_slice);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_15ce3046b2 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_15ce3046b2;


architecture behavior of relational_15ce3046b2 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_22_3_rel <= a_1_31 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub_wlan_phy_tx_pmd;
architecture behavior of xladdsub_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_60fd3b5996582b7a
    port (
          a: in std_logic_vector(9 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(9 - 1 downto 0)
    );
  end component;
  component addsb_11_0_d5bf78f2384e976c
    port (
          a: in std_logic_vector(10 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(10 - 1 downto 0)
    );
  end component;
  component addsb_11_0_8942e2ad5d8d4897
    port (
          a: in std_logic_vector(9 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(9 - 1 downto 0)
    );
  end component;
  component addsb_11_0_5c670787eb4ba225
    port (
          a: in std_logic_vector(3 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(3 - 1 downto 0)
    );
  end component;
  component addsb_11_0_a52ead9b8a3c1e76
    port (
          a: in std_logic_vector(9 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(9 - 1 downto 0)
    );
  end component;
  component addsb_11_0_7cf14debcedb76ce
    port (
          a: in std_logic_vector(13 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(13 - 1 downto 0)
    );
  end component;
  component addsb_11_0_73986f767e994888
    port (
          a: in std_logic_vector(10 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(10 - 1 downto 0)
    );
  end component;
  component addsb_11_0_7925f33378f00f6a
    port (
          a: in std_logic_vector(3 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(3 - 1 downto 0)
    );
  end component;
  component addsb_11_0_f66fe30ee2d0a6f0
    port (
          a: in std_logic_vector(17 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(17 - 1 downto 0)
    );
  end component;
  component addsb_11_0_6695c8a33176d3c2
    port (
          a: in std_logic_vector(18 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(18 - 1 downto 0)
    );
  end component;
  component addsb_11_0_2fe7f24afe1bc972
    port (
          a: in std_logic_vector(5 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(5 - 1 downto 0)
    );
  end component;
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_60fd3b5996582b7a")) generate
    core_instance0: addsb_11_0_60fd3b5996582b7a
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp1: if ((core_name0 = "addsb_11_0_d5bf78f2384e976c")) generate
    core_instance1: addsb_11_0_d5bf78f2384e976c
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_8942e2ad5d8d4897")) generate
    core_instance2: addsb_11_0_8942e2ad5d8d4897
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp3: if ((core_name0 = "addsb_11_0_5c670787eb4ba225")) generate
    core_instance3: addsb_11_0_5c670787eb4ba225
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp5: if ((core_name0 = "addsb_11_0_a52ead9b8a3c1e76")) generate
    core_instance5: addsb_11_0_a52ead9b8a3c1e76
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp6: if ((core_name0 = "addsb_11_0_7cf14debcedb76ce")) generate
    core_instance6: addsb_11_0_7cf14debcedb76ce
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp7: if ((core_name0 = "addsb_11_0_73986f767e994888")) generate
    core_instance7: addsb_11_0_73986f767e994888
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp8: if ((core_name0 = "addsb_11_0_7925f33378f00f6a")) generate
    core_instance8: addsb_11_0_7925f33378f00f6a
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp9: if ((core_name0 = "addsb_11_0_f66fe30ee2d0a6f0")) generate
    core_instance9: addsb_11_0_f66fe30ee2d0a6f0
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp10: if ((core_name0 = "addsb_11_0_6695c8a33176d3c2")) generate
    core_instance10: addsb_11_0_6695c8a33176d3c2
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp11: if ((core_name0 = "addsb_11_0_2fe7f24afe1bc972")) generate
    core_instance11: addsb_11_0_2fe7f24afe1bc972
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_305a9068e6 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_305a9068e6;


architecture behavior of relational_305a9068e6 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal cast_22_12: unsigned((9 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_12 <= u2u_cast(a_1_31, 0, 9, 0);
  result_22_3_rel <= cast_22_12 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a369e00c6b is
  port (
    in0 : in std_logic_vector((16 - 1) downto 0);
    in1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a369e00c6b;


architecture behavior of concat_a369e00c6b is
  signal in0_1_23: unsigned((16 - 1) downto 0);
  signal in1_1_27: unsigned((16 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_7025463ea8 is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_7025463ea8;


architecture behavior of reinterpret_7025463ea8 is
  signal input_port_1_40: signed((16 - 1) downto 0);
  signal output_port_5_5_force: unsigned((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_151459306d is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_151459306d;


architecture behavior of reinterpret_151459306d is
  signal input_port_1_40: unsigned((16 - 1) downto 0);
  signal output_port_5_5_force: signed((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlslice is
    generic (
        new_msb      : integer := 9;
        new_lsb      : integer := 1;
        x_width      : integer := 16;
        y_width      : integer := 8);
    port (
        x : in std_logic_vector (x_width-1 downto 0);
        y : out std_logic_vector (y_width-1 downto 0));
end xlslice;
architecture behavior of xlslice is
begin
    y <= x(new_msb downto new_lsb);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_37567836aa is
  port (
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_37567836aa;


architecture behavior of constant_37567836aa is
begin
  op <= "00000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xldpram_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    c_width_a: integer := 13;
    c_address_width_a: integer := 4;
    c_width_b: integer := 13;
    c_address_width_b: integer := 4;
    c_has_sinita: integer := 0;
    c_has_sinitb: integer := 0;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width_a - 1 downto 0);
    addra: in std_logic_vector(c_address_width_a - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    a_ce: in std_logic;
    a_clk: in std_logic;
    rsta: in std_logic_vector(0 downto 0) := (others => '0');
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    douta: out std_logic_vector(c_width_a - 1 downto 0);
    dinb: in std_logic_vector(c_width_b - 1 downto 0);
    addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
    web: in std_logic_vector(0 downto 0);
    b_ce: in std_logic;
    b_clk: in std_logic;
    rstb: in std_logic_vector(0 downto 0) := (others => '0');
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    doutb: out std_logic_vector(c_width_b - 1 downto 0)
  );
end xldpram_wlan_phy_tx_pmd;
architecture behavior of xldpram_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;

  signal core_addra: std_logic_vector(c_address_width_a - 1 downto 0);
  signal core_addrb: std_logic_vector(c_address_width_b - 1 downto 0);
  signal core_dina, core_douta, dly_douta:
    std_logic_vector(c_width_a - 1 downto 0);
  signal core_dinb, core_doutb, dly_doutb:
    std_logic_vector(c_width_b - 1 downto 0);
  signal core_wea, core_web: std_logic;
  signal core_a_ce, core_b_ce: std_logic;
  signal sinita, sinitb: std_logic;

  component bmg_72_e4abe4c74ea5aa02
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_e4abe4c74ea5aa02:
    component is true;
  attribute fpga_dont_touch of bmg_72_e4abe4c74ea5aa02:
    component is "true";
  attribute box_type of bmg_72_e4abe4c74ea5aa02:
    component  is "black_box";
  component bmg_72_30fab105208816ae
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_30fab105208816ae:
    component is true;
  attribute fpga_dont_touch of bmg_72_30fab105208816ae:
    component is "true";
  attribute box_type of bmg_72_30fab105208816ae:
    component  is "black_box";
begin
  core_addra <= addra;
  core_dina <= dina;
  douta <= dly_douta;
  core_wea <= wea(0);
  core_a_ce <= a_ce and ena(0);
  sinita <= rsta(0) and a_ce;

  core_addrb <= addrb;
  core_dinb <= dinb;
  doutb <= dly_doutb;
  core_web <= web(0);
  core_b_ce <= b_ce and enb(0);
  sinitb <= rstb(0) and b_ce;
  comp0: if ((core_name0 = "bmg_72_e4abe4c74ea5aa02")) generate
    core_instance0: bmg_72_e4abe4c74ea5aa02
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_30fab105208816ae")) generate
    core_instance1: bmg_72_30fab105208816ae
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  latency_test: if (latency > 2) generate
    regA: synth_reg
      generic map (
        width => c_width_a,
        latency => latency - 2
      )
      port map (
        i => core_douta,
        ce => core_a_ce,
        clr => '0',
        clk => a_clk,
        o => dly_douta
      );
    regB: synth_reg
      generic map (
        width => c_width_b,
        latency => latency - 2
      )
      port map (
        i => core_doutb,
        ce => core_b_ce,
        clr => '0',
        clk => b_clk,
        o => dly_doutb
      );
  end generate;
  latency1: if (latency <= 2) generate
    dly_douta <= core_douta;
    dly_doutb <= core_doutb;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfast_fourier_transform_886093b6a909385035fdd94c865209c9 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    event_data_in_channel_halt:out std_logic;
    event_data_out_channel_halt:out std_logic;
    event_fft_overflow:out std_logic;
    event_frame_started:out std_logic;
    event_status_channel_halt:out std_logic;
    event_tlast_missing:out std_logic;
    event_tlast_unexpected:out std_logic;
    m_axis_data_tdata_xk_im:out std_logic_vector(15 downto 0);
    m_axis_data_tdata_xk_re:out std_logic_vector(15 downto 0);
    m_axis_data_tlast:out std_logic;
    m_axis_data_tready:in std_logic;
    m_axis_data_tuser_ovflo:out std_logic_vector(0 downto 0);
    m_axis_data_tuser_xk_index:out std_logic_vector(5 downto 0);
    m_axis_data_tvalid:out std_logic;
    m_axis_status_tdata_ovflo:out std_logic_vector(0 downto 0);
    m_axis_status_tready:in std_logic;
    m_axis_status_tvalid:out std_logic;
    rst:in std_logic;
    s_axis_config_tdata_fwd_inv:in std_logic_vector(0 downto 0);
    s_axis_config_tdata_scale_sch:in std_logic_vector(5 downto 0);
    s_axis_config_tready:out std_logic;
    s_axis_config_tvalid:in std_logic;
    s_axis_data_tdata_xn_im:in std_logic_vector(15 downto 0);
    s_axis_data_tdata_xn_re:in std_logic_vector(15 downto 0);
    s_axis_data_tlast:in std_logic;
    s_axis_data_tready:out std_logic;
    s_axis_data_tvalid:in std_logic
  );
end xlfast_fourier_transform_886093b6a909385035fdd94c865209c9;


architecture behavior of xlfast_fourier_transform_886093b6a909385035fdd94c865209c9  is
  component xfft_v8_0_3683b4047ed128ab
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      aresetn:in std_logic;
      event_data_in_channel_halt:out std_logic;
      event_data_out_channel_halt:out std_logic;
      event_fft_overflow:out std_logic;
      event_frame_started:out std_logic;
      event_status_channel_halt:out std_logic;
      event_tlast_missing:out std_logic;
      event_tlast_unexpected:out std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tlast:out std_logic;
      m_axis_data_tready:in std_logic;
      m_axis_data_tuser:out std_logic_vector(15 downto 0);
      m_axis_data_tvalid:out std_logic;
      m_axis_status_tdata:out std_logic_vector(7 downto 0);
      m_axis_status_tready:in std_logic;
      m_axis_status_tvalid:out std_logic;
      s_axis_config_tdata:in std_logic_vector(7 downto 0);
      s_axis_config_tready:out std_logic;
      s_axis_config_tvalid:in std_logic;
      s_axis_data_tdata:in std_logic_vector(31 downto 0);
      s_axis_data_tlast:in std_logic;
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal aresetn_net: std_logic := '0';
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(15 downto 0) := (others=>'0');
signal m_axis_status_tdata_net: std_logic_vector(7 downto 0) := (others=>'0');
signal s_axis_config_tdata_net: std_logic_vector(7 downto 0) := (others=>'0');
signal s_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  aresetn_net <= rst or (not ce);
  m_axis_data_tdata_xk_im <= m_axis_data_tdata_net(31 downto 16);
  m_axis_data_tdata_xk_re <= m_axis_data_tdata_net(15 downto 0);
  m_axis_data_tuser_ovflo <= m_axis_data_tuser_net(8 downto 8);
  m_axis_data_tuser_xk_index <= m_axis_data_tuser_net(5 downto 0);
  m_axis_status_tdata_ovflo <= m_axis_status_tdata_net(0 downto 0);
  s_axis_config_tdata_net(6 downto 1) <= s_axis_config_tdata_scale_sch;
  s_axis_config_tdata_net(0 downto 0) <= s_axis_config_tdata_fwd_inv;
  s_axis_data_tdata_net(31 downto 16) <= s_axis_data_tdata_xn_im;
  s_axis_data_tdata_net(15 downto 0) <= s_axis_data_tdata_xn_re;
  xfft_v8_0_3683b4047ed128ab_instance : xfft_v8_0_3683b4047ed128ab
    port map(
      aclk=>clk,
      aclken=>ce,
      aresetn=>aresetn_net,
      event_data_in_channel_halt=>event_data_in_channel_halt,
      event_data_out_channel_halt=>event_data_out_channel_halt,
      event_fft_overflow=>event_fft_overflow,
      event_frame_started=>event_frame_started,
      event_status_channel_halt=>event_status_channel_halt,
      event_tlast_missing=>event_tlast_missing,
      event_tlast_unexpected=>event_tlast_unexpected,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tlast=>m_axis_data_tlast,
      m_axis_data_tready=>m_axis_data_tready,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid,
      m_axis_status_tdata=>m_axis_status_tdata_net,
      m_axis_status_tready=>m_axis_status_tready,
      m_axis_status_tvalid=>m_axis_status_tvalid,
      s_axis_config_tdata=>s_axis_config_tdata_net,
      s_axis_config_tready=>s_axis_config_tready,
      s_axis_config_tvalid=>s_axis_config_tvalid,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tlast=>s_axis_data_tlast,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>s_axis_data_tvalid
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.conv_pkg.all;
entity xlaxififogen_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    tdata_width: integer := -1;
    tdest_width: integer := -1;
    tstrb_width: integer := -1;
    tkeep_width: integer := -1;
    tid_width: integer := -1;
    tuser_width: integer := -1;
    has_aresetn: integer := -1;
    depth_bits: integer :=-1
  );
  port (
      s_aclk: in std_logic;
      ce: in std_logic;
      aresetn: in std_logic;
s_axis_tdata: in std_logic_vector(tdata_width - 1 downto 0):= (others => '0');
s_axis_tdest: in std_logic_vector(tdest_width - 1 downto 0):= (others => '0');
s_axis_tstrb: in std_logic_vector(tstrb_width - 1 downto 0):= (others => '0');
s_axis_tkeep: in std_logic_vector(tkeep_width - 1 downto 0):= (others => '0');
s_axis_tlast: in std_logic := '0';
s_axis_tid  : in std_logic_vector(tid_width - 1 downto 0):= (others => '0');
s_axis_tuser: in std_logic_vector(tuser_width - 1 downto 0):= (others => '0');
m_axis_tdata: out std_logic_vector(tdata_width - 1 downto 0);
m_axis_tdest: out std_logic_vector(tdest_width - 1 downto 0);
m_axis_tstrb: out std_logic_vector(tstrb_width - 1 downto 0);
m_axis_tkeep: out std_logic_vector(tkeep_width - 1 downto 0);
m_axis_tlast: out std_logic;
m_axis_tid  : out std_logic_vector(tid_width - 1 downto 0);
m_axis_tuser: out std_logic_vector(tuser_width - 1 downto 0);
      axis_underflow: out std_logic;
      axis_overflow: out std_logic;
      axis_data_count: out std_logic_vector( depth_bits - 1 downto 0);
      axis_prog_full_thresh: in std_logic_vector( depth_bits - 2 downto 0):= (others => '0');
      axis_prog_empty_thresh: in std_logic_vector(depth_bits - 2 downto 0):= (others => '0');

      s_axis_tvalid: in std_logic;
      s_axis_tready: out std_logic;
      m_axis_tready: in std_logic;
      m_axis_tvalid: out std_logic
  );
end xlaxififogen_wlan_phy_tx_pmd;
architecture behavior of xlaxififogen_wlan_phy_tx_pmd is
  component axififo_fg92_83e0abc99b742965
    port (
      s_aclk: in std_logic;
      s_aresetn: in std_logic;
      axis_data_count: out std_logic_vector( depth_bits - 1  downto 0);
      s_axis_tdata: in std_logic_vector(tdata_width - 1 downto 0);
      s_axis_tlast: in std_logic;
      s_axis_tuser: in std_logic_vector(tuser_width - 1 downto 0);
      s_axis_tvalid: in std_logic;
      s_axis_tready: out std_logic;
      m_axis_tdata: out std_logic_vector(tdata_width - 1 downto 0);
      m_axis_tlast: out std_logic;
      m_axis_tuser: out std_logic_vector(tuser_width - 1 downto 0);
      m_axis_tvalid: out std_logic;
      m_axis_tready: in std_logic

    );
  end component;

  attribute syn_black_box of axififo_fg92_83e0abc99b742965:
    component is true;
  attribute fpga_dont_touch of axififo_fg92_83e0abc99b742965:
    component is "true";
  attribute box_type of axififo_fg92_83e0abc99b742965:
    component  is "black_box";
  signal srst: std_logic:= '0';
  signal reset_gen1: std_logic  := '0';
  signal reset_gen_d1: std_logic        := '0';
  signal reset_gen_d2: std_logic := '0';
begin
  comp0: if ((core_name0 = "axififo_fg92_83e0abc99b742965")) generate
    core_instance0: axififo_fg92_83e0abc99b742965
      port map (
        s_aclk => s_aclk,
        s_aresetn => srst,
        axis_data_count => axis_data_count,
        s_axis_tdata => s_axis_tdata,
        s_axis_tlast => s_axis_tlast,
        s_axis_tuser => s_axis_tuser,
        s_axis_tvalid => s_axis_tvalid,
        s_axis_tready => s_axis_tready,
        m_axis_tdata => m_axis_tdata,
        m_axis_tlast => m_axis_tlast,
        m_axis_tuser => m_axis_tuser,
        m_axis_tvalid => m_axis_tvalid,
        m_axis_tready => m_axis_tready

      );
  end generate;
        srst <= reset_gen_d2 when (has_aresetn = 0)
                else not ( (not aresetn) and ce );
 process(s_aclk)
 begin
         if(s_aclk'event AND s_aclk = '1') then
                         reset_gen1 <= '1';
                         reset_gen_d1 <= reset_gen1;
                         reset_gen_d2 <= reset_gen_d1;
        end if;
 end process;

end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_35690eb8ec is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((16 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_35690eb8ec;


architecture behavior of mux_35690eb8ec is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((16 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((16 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= cast(d1_1_27, 11, 16, 15, xlSigned);
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_d99e59b6d4 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_d99e59b6d4;


architecture behavior of mux_d99e59b6d4 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic;
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= std_logic_to_vector(unregy_join_6_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_42c705c90b is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_42c705c90b;


architecture behavior of mux_42c705c90b is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_91ce9c6dac is
  port (
    in0 : in std_logic_vector((5 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((2 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_91ce9c6dac;


architecture behavior of concat_91ce9c6dac is
  signal in0_1_23: unsigned((5 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((2 - 1) downto 0);
  signal in4_1_39: boolean;
  signal in5_1_43: boolean;
  signal in6_1_47: boolean;
  signal in7_1_51: boolean;
  signal in8_1_55: boolean;
  signal y_2_1_concat: unsigned((18 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= ((in4) = "1");
  in5_1_43 <= ((in5) = "1");
  in6_1_47 <= ((in6) = "1");
  in7_1_51 <= ((in7) = "1");
  in8_1_55 <= ((in8) = "1");
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & boolean_to_vector(in4_1_39) & boolean_to_vector(in5_1_43) & boolean_to_vector(in6_1_47) & boolean_to_vector(in7_1_51) & boolean_to_vector(in8_1_55));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_ef0e2e5fc6 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_ef0e2e5fc6;


architecture behavior of constant_ef0e2e5fc6 is
begin
  op <= "10000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_469094441c is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_469094441c;


architecture behavior of constant_469094441c is
begin
  op <= "100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cda50df78a is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cda50df78a;


architecture behavior of constant_cda50df78a is
begin
  op <= "00";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_3a9a3daeb9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_3a9a3daeb9;


architecture behavior of constant_3a9a3daeb9 is
begin
  op <= "11";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fe72737ca0 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fe72737ca0;


architecture behavior of constant_fe72737ca0 is
begin
  op <= "00000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8ddc079e9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8ddc079e9;


architecture behavior of constant_e8ddc079e9 is
begin
  op <= "10";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4e64dfaf34 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4e64dfaf34;


architecture behavior of constant_4e64dfaf34 is
begin
  op <= "101";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_2a63ac73aa is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_2a63ac73aa;


architecture behavior of mux_2a63ac73aa is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((2 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_1d0997f32b is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_1d0997f32b;


architecture behavior of relational_1d0997f32b is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_12_17: unsigned((10 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_0f9b7ba263 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_0f9b7ba263;


architecture behavior of relational_0f9b7ba263 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_20_17: unsigned((10 - 1) downto 0);
  signal result_20_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_20_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_20_3_rel <= a_1_31 <= cast_20_17;
  op <= boolean_to_vector(result_20_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_3c449faea2 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_3c449faea2;


architecture behavior of relational_3c449faea2 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_22_17: unsigned((10 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_22_3_rel <= a_1_31 >= cast_22_17;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_7907e32f0f is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_7907e32f0f;


architecture behavior of relational_7907e32f0f is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_22_17: unsigned((10 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_22_3_rel <= a_1_31 >= cast_22_17;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9108cf519a is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9108cf519a;


architecture behavior of relational_9108cf519a is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_12_17: unsigned((10 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5b4e5df320 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5b4e5df320;


architecture behavior of relational_5b4e5df320 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_12_17: unsigned((10 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6158158994 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6158158994;


architecture behavior of relational_6158158994 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal cast_22_17: unsigned((10 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_17 <= u2u_cast(b_1_34, 0, 10, 0);
  result_22_3_rel <= a_1_31 >= cast_22_17;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b8fb990c43 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b8fb990c43;


architecture behavior of constant_b8fb990c43 is
begin
  op <= "10110100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_a6d07705dd is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_a6d07705dd;


architecture behavior of logical_a6d07705dd is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal d3_1_33: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  d3_1_33 <= d3(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27 or d2_1_30 or d3_1_33;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_954ee29728 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_954ee29728;


architecture behavior of logical_954ee29728 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27 and d2_1_30;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_ecce2f20df is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_ecce2f20df;


architecture behavior of relational_ecce2f20df is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_16_16: unsigned((10 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_16_16 <= u2u_cast(b_1_34, 0, 10, 0);
  result_16_3_rel <= a_1_31 < cast_16_16;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2d417722ee is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2d417722ee;


architecture behavior of relational_2d417722ee is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_20_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_20_3_rel <= a_1_31 <= b_1_34;
  op <= boolean_to_vector(result_20_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_899cf9b568 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_899cf9b568;


architecture behavior of logical_899cf9b568 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal d3_1_33: std_logic_vector((1 - 1) downto 0);
  signal d4_1_36: std_logic_vector((1 - 1) downto 0);
  signal en_1_39: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (1 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    0 => "0");
  signal latency_pipe_5_26_front_din: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_back: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_shift_join_7_1: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_shift_join_7_1_en: std_logic;
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  en_1_39 <= en(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(0);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  fully_2_1_bit <= d0_1_24 xor d1_1_27 xor d2_1_30 xor d3_1_33 xor d4_1_36;
  proc_if_7_1: process (en_1_39, fully_2_1_bit)
  is
  begin
    if en_1_39 = '1' then
      latency_pipe_shift_join_7_1_en <= '1';
    else 
      latency_pipe_shift_join_7_1_en <= '0';
    end if;
    latency_pipe_shift_join_7_1 <= fully_2_1_bit;
  end process proc_if_7_1;
  latency_pipe_5_26_front_din <= latency_pipe_shift_join_7_1;
  latency_pipe_5_26_push_front_pop_back_en <= latency_pipe_shift_join_7_1_en;
  y <= latency_pipe_5_26_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_706b9eb7ce is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_706b9eb7ce;


architecture behavior of relational_706b9eb7ce is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_12_17: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 3, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_bc74ae1a6c is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_bc74ae1a6c;


architecture behavior of constant_bc74ae1a6c is
begin
  op <= "11000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_02d5ef99fc is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((10 - 1) downto 0);
    d1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_02d5ef99fc;


architecture behavior of mux_02d5ef99fc is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((10 - 1) downto 0);
  signal d1_1_27: std_logic_vector((5 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((10 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= cast(d1_1_27, 0, 10, 0, xlUnsigned);
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_1813613113 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_1813613113;


architecture behavior of relational_1813613113 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd8727242d is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd8727242d;


architecture behavior of constant_fd8727242d is
begin
  op <= "011100000111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c09b53cba3 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c09b53cba3;


architecture behavior of constant_c09b53cba3 is
begin
  op <= "100011111001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_41d1fb8f4c is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_41d1fb8f4c;


architecture behavior of constant_41d1fb8f4c is
begin
  op <= "110110101000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_aec943c743 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_aec943c743;


architecture behavior of constant_aec943c743 is
begin
  op <= "001001011000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_192c5da026 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    d3 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_192c5da026;


architecture behavior of mux_192c5da026 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal d3_1_33: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9127ce6619 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9127ce6619;


architecture behavior of constant_9127ce6619 is
begin
  op <= "011111111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_50239c0b0e is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_50239c0b0e;


architecture behavior of constant_50239c0b0e is
begin
  op <= "101001001001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1971ed2879 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1971ed2879;


architecture behavior of constant_1971ed2879 is
begin
  op <= "110010010010";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_93635891b9 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_93635891b9;


architecture behavior of constant_93635891b9 is
begin
  op <= "001101101110";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e054d850c5 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e054d850c5;


architecture behavior of constant_e054d850c5 is
begin
  op <= "100000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9fcec64691 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9fcec64691;


architecture behavior of constant_9fcec64691 is
begin
  op <= "111011011011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8da791e271 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8da791e271;


architecture behavior of constant_8da791e271 is
begin
  op <= "000100100101";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c3ad5f20a9 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c3ad5f20a9;


architecture behavior of constant_c3ad5f20a9 is
begin
  op <= "010110110111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f3bb14635d is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    d3 : in std_logic_vector((12 - 1) downto 0);
    d4 : in std_logic_vector((12 - 1) downto 0);
    d5 : in std_logic_vector((12 - 1) downto 0);
    d6 : in std_logic_vector((12 - 1) downto 0);
    d7 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f3bb14635d;


architecture behavior of mux_f3bb14635d is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal d3_1_33: std_logic_vector((12 - 1) downto 0);
  signal d4_1_36: std_logic_vector((12 - 1) downto 0);
  signal d5_1_39: std_logic_vector((12 - 1) downto 0);
  signal d6_1_42: std_logic_vector((12 - 1) downto 0);
  signal d7_1_45: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7e4d1a10e6 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7e4d1a10e6;


architecture behavior of constant_7e4d1a10e6 is
begin
  op <= "100010011000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_afc893bf70 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_afc893bf70;


architecture behavior of constant_afc893bf70 is
begin
  op <= "011101101000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd28b32bf8 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd28b32bf8;


architecture behavior of constant_fd28b32bf8 is
begin
  op <= "000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_c3e1ddb86e is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_c3e1ddb86e;


architecture behavior of mux_c3e1ddb86e is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4de2214a42 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4de2214a42;


architecture behavior of mux_4de2214a42 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7b07120b87 is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7b07120b87;


architecture behavior of constant_7b07120b87 is
begin
  op <= "1000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_3797c120ed is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((7 - 1) downto 0);
    d1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_3797c120ed;


architecture behavior of mux_3797c120ed is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((7 - 1) downto 0);
  signal d1_1_27: std_logic_vector((7 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((7 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_23065a6aa3 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_23065a6aa3;


architecture behavior of relational_23065a6aa3 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1f05b15a2d is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1f05b15a2d;


architecture behavior of constant_1f05b15a2d is
begin
  op <= "010101";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_330e503d71 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_330e503d71;


architecture behavior of constant_330e503d71 is
begin
  op <= "000111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_173d83e4a7 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_173d83e4a7;


architecture behavior of constant_173d83e4a7 is
begin
  op <= "111001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8207020ee3 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8207020ee3;


architecture behavior of constant_8207020ee3 is
begin
  op <= "101011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_cdffdf53c9 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_cdffdf53c9;


architecture behavior of mux_cdffdf53c9 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal d3_1_33: std_logic;
  signal unregy_join_6_1: std_logic;
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  d3_1_33 <= d3(0);
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= std_logic_to_vector(unregy_join_6_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_931d61fb72 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_931d61fb72;


architecture behavior of relational_931d61fb72 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlpassthrough is
    generic (
        din_width    : integer := 16;
        dout_width   : integer := 16
        );
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlpassthrough;
architecture passthrough_arch of xlpassthrough is
begin
  dout <= din;
end passthrough_arch;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_e77c53f8bd is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_e77c53f8bd;


architecture behavior of logical_e77c53f8bd is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_47932db5b1 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_47932db5b1;


architecture behavior of relational_47932db5b1 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_1834ac00b4 is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_1834ac00b4;


architecture behavior of relational_1834ac00b4 is
  signal a_1_31: signed((9 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal cast_12_17: signed((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_signed(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2s_cast(b_1_34, 0, 9, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_32afb77cd2 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_32afb77cd2;


architecture behavior of concat_32afb77cd2 is
  signal in0_1_23: boolean;
  signal in1_1_27: boolean;
  signal y_2_1_concat: unsigned((2 - 1) downto 0);
begin
  in0_1_23 <= ((in0) = "1");
  in1_1_27 <= ((in1) = "1");
  y_2_1_concat <= std_logic_vector_to_unsigned(boolean_to_vector(in0_1_23) & boolean_to_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cb767c7ef2 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cb767c7ef2;


architecture behavior of constant_cb767c7ef2 is
begin
  op <= "101011000011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_d6a72b7a3b is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_d6a72b7a3b;


architecture behavior of constant_d6a72b7a3b is
begin
  op <= "010100111101";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_33c9a0c803 is
  port (
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_33c9a0c803;


architecture behavior of logical_33c9a0c803 is
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((2 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_e5a9964709 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_e5a9964709;


architecture behavior of mux_e5a9964709 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c0ce4ae10c is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c0ce4ae10c;


architecture behavior of constant_c0ce4ae10c is
begin
  op <= "1011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_5c1626e05e is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_5c1626e05e;


architecture behavior of constant_5c1626e05e is
begin
  op <= "1010";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1e60cf48bc is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((3 - 1) downto 0);
    d1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1e60cf48bc;


architecture behavior of mux_1e60cf48bc is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((3 - 1) downto 0);
  signal d1_1_27: std_logic_vector((4 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((4 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 4, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_102f86419c is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((4 - 1) downto 0);
    d1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_102f86419c;


architecture behavior of mux_102f86419c is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((4 - 1) downto 0);
  signal d1_1_27: std_logic_vector((3 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((4 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= cast(d1_1_27, 0, 4, 0, xlUnsigned);
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_b218b04ee6 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_b218b04ee6;


architecture behavior of relational_b218b04ee6 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal cast_20_17: unsigned((12 - 1) downto 0);
  signal result_20_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_20_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_20_3_rel <= a_1_31 <= cast_20_17;
  op <= boolean_to_vector(result_20_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c5804edea5 is
  port (
    in0 : in std_logic_vector((16 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    in2 : in std_logic_vector((9 - 1) downto 0);
    in3 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c5804edea5;


architecture behavior of concat_c5804edea5 is
  signal in0_1_23: unsigned((16 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal in2_1_31: unsigned((9 - 1) downto 0);
  signal in3_1_35: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_822933f89b is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_822933f89b;


architecture behavior of constant_822933f89b is
begin
  op <= "000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9f5572ba51 is
  port (
    op : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9f5572ba51;


architecture behavior of constant_9f5572ba51 is
begin
  op <= "0000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c4c603edf2 is
  port (
    op : out std_logic_vector((64 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c4c603edf2;


architecture behavior of constant_c4c603edf2 is
begin
  op <= "0000000000000000000000000000000000000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_91ef1678ca is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_91ef1678ca;


architecture behavior of constant_91ef1678ca is
begin
  op <= "00000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_c762ea476a is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    d2 : in std_logic_vector((8 - 1) downto 0);
    d3 : in std_logic_vector((8 - 1) downto 0);
    d4 : in std_logic_vector((8 - 1) downto 0);
    d5 : in std_logic_vector((8 - 1) downto 0);
    d6 : in std_logic_vector((8 - 1) downto 0);
    d7 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_c762ea476a;


architecture behavior of mux_c762ea476a is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal d2_1_30: std_logic_vector((8 - 1) downto 0);
  signal d3_1_33: std_logic_vector((8 - 1) downto 0);
  signal d4_1_36: std_logic_vector((8 - 1) downto 0);
  signal d5_1_39: std_logic_vector((8 - 1) downto 0);
  signal d6_1_42: std_logic_vector((8 - 1) downto 0);
  signal d7_1_45: std_logic_vector((8 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((8 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_b0082e75ff is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    d5 : in std_logic_vector((1 - 1) downto 0);
    d6 : in std_logic_vector((1 - 1) downto 0);
    d7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_b0082e75ff;


architecture behavior of mux_b0082e75ff is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal d3_1_33: std_logic_vector((1 - 1) downto 0);
  signal d4_1_36: std_logic_vector((1 - 1) downto 0);
  signal d5_1_39: std_logic_vector((1 - 1) downto 0);
  signal d6_1_42: std_logic_vector((1 - 1) downto 0);
  signal d7_1_45: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((1 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_998e20a1ca is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    d2 : in std_logic_vector((8 - 1) downto 0);
    d3 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_998e20a1ca;


architecture behavior of mux_998e20a1ca is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal d2_1_30: std_logic_vector((8 - 1) downto 0);
  signal d3_1_33: std_logic_vector((8 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((8 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_387191112d is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_387191112d;


architecture behavior of mux_387191112d is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((8 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7673b9b993 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7673b9b993;


architecture behavior of concat_7673b9b993 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a1e126f11c is
  port (
    in0 : in std_logic_vector((8 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    in2 : in std_logic_vector((8 - 1) downto 0);
    in3 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a1e126f11c;


architecture behavior of concat_a1e126f11c is
  signal in0_1_23: unsigned((8 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal in2_1_31: unsigned((8 - 1) downto 0);
  signal in3_1_35: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c048fbe4a5 is
  port (
    in0 : in std_logic_vector((24 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c048fbe4a5;


architecture behavior of concat_c048fbe4a5 is
  signal in0_1_23: unsigned((24 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_6a3d3dd4e5 is
  port (
    ip : in std_logic_vector((32 - 1) downto 0);
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_6a3d3dd4e5;


architecture behavior of inverter_6a3d3dd4e5 is
  signal ip_1_26: unsigned((32 - 1) downto 0);
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of unsigned((32 - 1) downto 0);
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => "00000000000000000000000000000000");
  signal op_mem_22_20_front_din: unsigned((32 - 1) downto 0);
  signal op_mem_22_20_back: unsigned((32 - 1) downto 0);
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: unsigned((32 - 1) downto 0);
begin
  ip_1_26 <= std_logic_vector_to_unsigned(ip);
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= std_logic_vector_to_unsigned(not unsigned_to_std_logic_vector(ip_1_26));
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_59f8d33339 is
  port (
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_59f8d33339;


architecture behavior of logical_59f8d33339 is
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((8 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_b23aa74086 is
  port (
    d0 : in std_logic_vector((32 - 1) downto 0);
    d1 : in std_logic_vector((32 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_b23aa74086;


architecture behavior of logical_b23aa74086 is
  signal d0_1_24: std_logic_vector((32 - 1) downto 0);
  signal d1_1_27: std_logic_vector((32 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((32 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_28e8664d0c is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_28e8664d0c;


architecture behavior of relational_28e8664d0c is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal cast_22_17: unsigned((12 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_22_3_rel <= a_1_31 >= cast_22_17;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_ae4e737ca0 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_ae4e737ca0;


architecture behavior of relational_ae4e737ca0 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_22_17: unsigned((12 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_22_3_rel <= a_1_31 >= cast_22_17;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0f59f02ba5 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0f59f02ba5;


architecture behavior of constant_0f59f02ba5 is
begin
  op <= "011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a629aefb53 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a629aefb53;


architecture behavior of constant_a629aefb53 is
begin
  op <= "1001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_263f209841 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_263f209841;


architecture behavior of constant_263f209841 is
begin
  op <= "110";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1f5cc32f1e is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1f5cc32f1e;


architecture behavior of constant_1f5cc32f1e is
begin
  op <= "010";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8038205d89 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8038205d89;


architecture behavior of constant_8038205d89 is
begin
  op <= "0011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_82200c2969 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_82200c2969;


architecture behavior of relational_82200c2969 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: signed((18 - 1) downto 0);
  signal cast_22_12: signed((18 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_signed(b);
  cast_22_12 <= u2s_cast(a_1_31, 0, 18, 0);
  result_22_3_rel <= cast_22_12 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_31ab9f25e5 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_31ab9f25e5;


architecture behavior of relational_31ab9f25e5 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal cast_16_16: unsigned((12 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_16_16 <= u2u_cast(b_1_34, 0, 12, 0);
  result_16_3_rel <= a_1_31 < cast_16_16;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_61c9d3f3fc is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((17 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_61c9d3f3fc;


architecture behavior of relational_61c9d3f3fc is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((17 - 1) downto 0);
  signal cast_22_12: unsigned((17 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_12 <= u2u_cast(a_1_31, 0, 17, 0);
  result_22_3_rel <= cast_22_12 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_ab46f67027 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((17 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_ab46f67027;


architecture behavior of relational_ab46f67027 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((17 - 1) downto 0);
  signal cast_12_12: unsigned((17 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_12 <= u2u_cast(a_1_31, 0, 17, 0);
  result_12_3_rel <= cast_12_12 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6c709b1b0c is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6c709b1b0c;


architecture behavior of relational_6c709b1b0c is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0c7cd7a34 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0c7cd7a34;


architecture behavior of concat_a0c7cd7a34 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_9d76333483 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_9d76333483;


architecture behavior of logical_9d76333483 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_1a070f1f35 is
  port (
    in0 : in std_logic_vector((4 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_1a070f1f35;


architecture behavior of concat_1a070f1f35 is
  signal in0_1_23: unsigned((4 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_bfd5ba0f50 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_bfd5ba0f50;


architecture behavior of constant_bfd5ba0f50 is
begin
  op <= "0110";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_4a6def08e4 is
  port (
    ip : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_4a6def08e4;


architecture behavior of inverter_4a6def08e4 is
  signal ip_1_26: unsigned((8 - 1) downto 0);
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of unsigned((8 - 1) downto 0);
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => "00000000");
  signal op_mem_22_20_front_din: unsigned((8 - 1) downto 0);
  signal op_mem_22_20_back: unsigned((8 - 1) downto 0);
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: unsigned((8 - 1) downto 0);
begin
  ip_1_26 <= std_logic_vector_to_unsigned(ip);
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= std_logic_vector_to_unsigned(not unsigned_to_std_logic_vector(ip_1_26));
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_dc245eb1d2 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_dc245eb1d2;


architecture behavior of concat_dc245eb1d2 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7ea0f2fff7 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7ea0f2fff7;


architecture behavior of constant_7ea0f2fff7 is
begin
  op <= "000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_8e53793314 is
  port (
    in0 : in std_logic_vector((8 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_8e53793314;


architecture behavior of concat_8e53793314 is
  signal in0_1_23: unsigned((8 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((16 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_0ee569a826 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_0ee569a826;


architecture behavior of logical_0ee569a826 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal d3_1_33: std_logic;
  signal d4_1_36: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  d3_1_33 <= d3(0);
  d4_1_36 <= d4(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27 or d2_1_30 or d3_1_33 or d4_1_36;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2a3f3bef9d is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2a3f3bef9d;


architecture behavior of relational_2a3f3bef9d is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_14_17: unsigned((2 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_14_17 <= u2u_cast(b_1_34, 0, 2, 0);
  result_14_3_rel <= a_1_31 /= cast_14_17;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ac785d9b37 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ac785d9b37;


architecture behavior of concat_ac785d9b37 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1d6ad1c713 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1d6ad1c713;


architecture behavior of constant_1d6ad1c713 is
begin
  op <= "111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1a631d900c is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1a631d900c;


architecture behavior of constant_1a631d900c is
begin
  op <= "0011111";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_wlan_phy_tx_pmd ;
architecture behavior of xlsprom_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_ce, sinit: std_logic;
  component bmg_72_d44417b0abe027bf
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_d44417b0abe027bf:
    component is true;
  attribute fpga_dont_touch of bmg_72_d44417b0abe027bf:
    component is "true";
  attribute box_type of bmg_72_d44417b0abe027bf:
    component  is "black_box";
  component bmg_72_8bdf24f02e925a98
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_8bdf24f02e925a98:
    component is true;
  attribute fpga_dont_touch of bmg_72_8bdf24f02e925a98:
    component is "true";
  attribute box_type of bmg_72_8bdf24f02e925a98:
    component  is "black_box";
begin
  core_addr <= addr;
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_d44417b0abe027bf")) generate
    core_instance0: bmg_72_d44417b0abe027bf
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp1: if ((core_name0 = "bmg_72_8bdf24f02e925a98")) generate
    core_instance1: bmg_72_8bdf24f02e925a98
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_1: if (latency <= 1) generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_c5ffb0182e is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_c5ffb0182e;


architecture behavior of relational_c5ffb0182e is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_18_16: unsigned((7 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_18_16 <= u2u_cast(b_1_34, 0, 7, 0);
  result_18_3_rel <= a_1_31 > cast_18_16;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_27dbff5dcf is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_27dbff5dcf;


architecture behavior of relational_27dbff5dcf is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_20_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_20_3_rel <= a_1_31 <= b_1_34;
  op <= boolean_to_vector(result_20_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_145086465d is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_145086465d;


architecture behavior of constant_145086465d is
begin
  op <= "1000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f1cd62c228 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    d2 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f1cd62c228;


architecture behavior of mux_f1cd62c228 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal d2_1_30: std_logic_vector((8 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((8 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_09ceb5d9bd is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_09ceb5d9bd;


architecture behavior of relational_09ceb5d9bd is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_12_17: unsigned((12 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_ae8b814968 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_ae8b814968;


architecture behavior of relational_ae8b814968 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_12_17: unsigned((12 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5321bc1192 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5321bc1192;


architecture behavior of relational_5321bc1192 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal cast_12_17: unsigned((12 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 12, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_1d9bdbb01e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    in2 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_1d9bdbb01e;


architecture behavior of concat_1d9bdbb01e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal in2_1_31: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a1c496ea88 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a1c496ea88;


architecture behavior of constant_a1c496ea88 is
begin
  op <= "001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_8a8a6c93e0 is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((3 - 1) downto 0);
    d1 : in std_logic_vector((3 - 1) downto 0);
    d2 : in std_logic_vector((3 - 1) downto 0);
    d3 : in std_logic_vector((3 - 1) downto 0);
    d4 : in std_logic_vector((3 - 1) downto 0);
    d5 : in std_logic_vector((3 - 1) downto 0);
    d6 : in std_logic_vector((3 - 1) downto 0);
    d7 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_8a8a6c93e0;


architecture behavior of mux_8a8a6c93e0 is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((3 - 1) downto 0);
  signal d1_1_27: std_logic_vector((3 - 1) downto 0);
  signal d2_1_30: std_logic_vector((3 - 1) downto 0);
  signal d3_1_33: std_logic_vector((3 - 1) downto 0);
  signal d4_1_36: std_logic_vector((3 - 1) downto 0);
  signal d5_1_39: std_logic_vector((3 - 1) downto 0);
  signal d6_1_42: std_logic_vector((3 - 1) downto 0);
  signal d7_1_45: std_logic_vector((3 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((3 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_9ac2bdb119 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    d5 : in std_logic_vector((1 - 1) downto 0);
    d6 : in std_logic_vector((1 - 1) downto 0);
    d7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_9ac2bdb119;


architecture behavior of logical_9ac2bdb119 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal d3_1_33: std_logic_vector((1 - 1) downto 0);
  signal d4_1_36: std_logic_vector((1 - 1) downto 0);
  signal d5_1_39: std_logic_vector((1 - 1) downto 0);
  signal d6_1_42: std_logic_vector((1 - 1) downto 0);
  signal d7_1_45: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  fully_2_1_bit <= d0_1_24 xor d1_1_27 xor d2_1_30 xor d3_1_33 xor d4_1_36 xor d5_1_39 xor d6_1_42 xor d7_1_45;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_604045dd09 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_604045dd09;


architecture behavior of logical_604045dd09 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  fully_2_1_bit <= d0_1_24 xor d1_1_27 xor d2_1_30;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_c49d820dc8 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_c49d820dc8;


architecture behavior of relational_c49d820dc8 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_14_17: unsigned((6 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_14_17 <= u2u_cast(b_1_34, 0, 6, 0);
  result_14_3_rel <= a_1_31 /= cast_14_17;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a7e2bb9e12 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a7e2bb9e12;


architecture behavior of constant_a7e2bb9e12 is
begin
  op <= "01";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_6cb8f0ce02 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_6cb8f0ce02;


architecture behavior of logical_6cb8f0ce02 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27 or d2_1_30;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_eb88ab7682 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((10 - 1) downto 0);
    d1 : in std_logic_vector((10 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_eb88ab7682;


architecture behavior of mux_eb88ab7682 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((10 - 1) downto 0);
  signal d1_1_27: std_logic_vector((10 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((10 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_a585e6d5ba is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_a585e6d5ba;


architecture behavior of mux_a585e6d5ba is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((16 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((16 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 16, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_938d99ac11 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_938d99ac11;


architecture behavior of logical_938d99ac11 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_13241d6573 is
  port (
    in0 : in std_logic_vector((6 - 1) downto 0);
    in1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_13241d6573;


architecture behavior of concat_13241d6573 is
  signal in0_1_23: unsigned((6 - 1) downto 0);
  signal in1_1_27: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_791081a00e is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((9 - 1) downto 0);
    d1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_791081a00e;


architecture behavior of mux_791081a00e is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((9 - 1) downto 0);
  signal d1_1_27: std_logic_vector((9 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((9 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity accum_3520344abf is
  port (
    b : in std_logic_vector((2 - 1) downto 0);
    rst : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end accum_3520344abf;


architecture behavior of accum_3520344abf is
  signal b_17_24: unsigned((2 - 1) downto 0);
  signal rst_17_27: boolean;
  signal en_17_32: boolean;
  signal accum_reg_41_23: unsigned((9 - 1) downto 0) := "000000000";
  signal accum_reg_41_23_rst: std_logic;
  signal accum_reg_41_23_en: std_logic;
  signal cast_51_42: unsigned((9 - 1) downto 0);
  signal accum_reg_join_47_1: unsigned((10 - 1) downto 0);
  signal accum_reg_join_47_1_en: std_logic;
  signal accum_reg_join_47_1_rst: std_logic;
begin
  b_17_24 <= std_logic_vector_to_unsigned(b);
  rst_17_27 <= ((rst) = "1");
  en_17_32 <= ((en) = "1");
  proc_accum_reg_41_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (accum_reg_41_23_rst = '1')) then
        accum_reg_41_23 <= "000000000";
      elsif ((ce = '1') and (accum_reg_41_23_en = '1')) then 
        accum_reg_41_23 <= accum_reg_41_23 + cast_51_42;
      end if;
    end if;
  end process proc_accum_reg_41_23;
  cast_51_42 <= u2u_cast(b_17_24, 0, 9, 0);
  proc_if_47_1: process (accum_reg_41_23, cast_51_42, en_17_32, rst_17_27)
  is
  begin
    if rst_17_27 then
      accum_reg_join_47_1_rst <= '1';
    elsif en_17_32 then
      accum_reg_join_47_1_rst <= '0';
    else 
      accum_reg_join_47_1_rst <= '0';
    end if;
    if en_17_32 then
      accum_reg_join_47_1_en <= '1';
    else 
      accum_reg_join_47_1_en <= '0';
    end if;
  end process proc_if_47_1;
  accum_reg_41_23_rst <= accum_reg_join_47_1_rst;
  accum_reg_41_23_en <= accum_reg_join_47_1_en;
  q <= unsigned_to_std_logic_vector(accum_reg_41_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2d0bbe9efa is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((2 - 1) downto 0);
    in2 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2d0bbe9efa;


architecture behavior of concat_2d0bbe9efa is
  signal in0_1_23: boolean;
  signal in1_1_27: unsigned((2 - 1) downto 0);
  signal in2_1_31: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= ((in0) = "1");
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(boolean_to_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd85eb7067 is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd85eb7067;


architecture behavior of constant_fd85eb7067 is
begin
  op <= "000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_194eb61c1b is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_194eb61c1b;


architecture behavior of relational_194eb61c1b is
  signal a_1_31: unsigned((1 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_12_12: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_12 <= u2u_cast(a_1_31, 0, 2, 0);
  result_12_3_rel <= cast_12_12 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_caa2b01eef is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_caa2b01eef;


architecture behavior of counter_caa2b01eef is
  signal rst_1_40: boolean;
  signal en_1_45: boolean;
  signal count_reg_20_23: unsigned((1 - 1) downto 0) := "0";
  signal count_reg_20_23_rst: std_logic;
  signal count_reg_20_23_en: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((2 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0";
      elsif ((ce = '1') and (count_reg_20_23_en = '1')) then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("1");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23, en_1_45)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    elsif en_1_45 then
      count_reg_join_44_1_rst <= '0';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    elsif en_1_45 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_78aa6a36ae is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    d2 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_78aa6a36ae;


architecture behavior of mux_78aa6a36ae is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal d2_1_30: std_logic_vector((2 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((2 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5f1eb17108 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5f1eb17108;


architecture behavior of relational_5f1eb17108 is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_f52e6abf76 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_f52e6abf76;


architecture behavior of relational_f52e6abf76 is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_12_17: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 2, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
entity xlcounter_limit_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned;
    cnt_63_48: integer:= 0;
    cnt_47_32: integer:= 0;
    cnt_31_16: integer:= 0;
    cnt_15_0: integer:= 0;
    count_limited: integer := 0
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_limit_wlan_phy_tx_pmd ;
architecture behavior of xlcounter_limit_wlan_phy_tx_pmd is
  signal high_cnt_to: std_logic_vector(31 downto 0);
  signal low_cnt_to: std_logic_vector(31 downto 0);
  signal cnt_to: std_logic_vector(63 downto 0);
  signal core_sinit, op_thresh0, core_ce: std_logic;
  signal rst_overrides_en: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
  -- synopsys translate_off
  signal real_op : real;
   -- synopsys translate_on
  function equals(op, cnt_to : std_logic_vector; width, arith : integer)
    return std_logic
  is
    variable signed_op, signed_cnt_to : signed (width - 1 downto 0);
    variable unsigned_op, unsigned_cnt_to : unsigned (width - 1 downto 0);
    variable result : std_logic;
  begin
    -- synopsys translate_off
    if ((is_XorU(op)) or (is_XorU(cnt_to)) ) then
      result := '0';
      return result;
    end if;
    -- synopsys translate_on
    if (op = cnt_to) then
      result := '1';
    else
      result := '0';
    end if;
    return result;
  end;
  component cntr_11_0_6454489cfe866515
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_6454489cfe866515:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_6454489cfe866515:
    component is "true";
  attribute box_type of cntr_11_0_6454489cfe866515:
    component  is "black_box";
  component cntr_11_0_bcc28bfecf25caff
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_bcc28bfecf25caff:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_bcc28bfecf25caff:
    component is "true";
  attribute box_type of cntr_11_0_bcc28bfecf25caff:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec : std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec : std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
begin
  -- synopsys translate_off
  -- synopsys translate_on
  cnt_to(63 downto 48) <= integer_to_std_logic_vector(cnt_63_48, 16, op_arith);
  cnt_to(47 downto 32) <= integer_to_std_logic_vector(cnt_47_32, 16, op_arith);
  cnt_to(31 downto 16) <= integer_to_std_logic_vector(cnt_31_16, 16, op_arith);
  cnt_to(15 downto 0) <= integer_to_std_logic_vector(cnt_15_0, 16, op_arith);
  op <= op_net;
  core_ce <= ce and en(0);
  rst_overrides_en <= rst(0) or en(0);
  limit : if (count_limited = 1) generate
    eq_cnt_to : process (op_net, cnt_to)
    begin
      op_thresh0 <= equals(op_net, cnt_to(op_width - 1 downto 0),
                     op_width, op_arith);
    end process;
    core_sinit <= (op_thresh0 or clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  no_limit : if (count_limited = 0) generate
    core_sinit <= (clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  comp0: if ((core_name0 = "cntr_11_0_6454489cfe866515")) generate
    core_instance0: cntr_11_0_6454489cfe866515
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_bcc28bfecf25caff")) generate
    core_instance1: cntr_11_0_bcc28bfecf25caff
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_8fc7f5539b is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_8fc7f5539b;


architecture behavior of relational_8fc7f5539b is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1a0db76efe is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    d2 : in std_logic_vector((2 - 1) downto 0);
    d3 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1a0db76efe;


architecture behavior of mux_1a0db76efe is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal d2_1_30: std_logic_vector((2 - 1) downto 0);
  signal d3_1_33: std_logic_vector((2 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((2 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.conv_pkg.all;
entity xlfifogen_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    data_width: integer := -1;
    data_count_width: integer := -1;
    percent_full_width: integer := -1;
    has_ae : integer := 0;
    has_af : integer := 0
  );
  port (
    din: in std_logic_vector(data_width - 1 downto 0);
    we: in std_logic;
    we_ce: in std_logic;
    re: in std_logic;
    re_ce: in std_logic;
    rst: in std_logic;
    en: in std_logic;
    ce: in std_logic;
    clk: in std_logic;
    empty: out std_logic;
    full: out std_logic;
    percent_full: out std_logic_vector(percent_full_width - 1 downto 0);
    dcount: out std_logic_vector(data_count_width - 1 downto 0);
    ae: out std_logic;
    af: out std_logic;
    dout: out std_logic_vector(data_width - 1 downto 0)
  );
end xlfifogen_wlan_phy_tx_pmd ;
architecture behavior of xlfifogen_wlan_phy_tx_pmd is
  component fifo_fg92_6a1156e8dc43a711
    port (
      clk: in std_logic;
      srst: in std_logic;
      din: in std_logic_vector(data_width - 1 downto 0);
      wr_en: in std_logic;
      rd_en: in std_logic;
      dout: out std_logic_vector(data_width - 1 downto 0);
      full: out std_logic;
      empty: out std_logic;
      data_count: out std_logic_vector(data_count_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of fifo_fg92_6a1156e8dc43a711:
    component is true;
  attribute fpga_dont_touch of fifo_fg92_6a1156e8dc43a711:
    component is "true";
  attribute box_type of fifo_fg92_6a1156e8dc43a711:
    component  is "black_box";
  signal rd_en: std_logic;
  signal wr_en: std_logic;
  signal srst: std_logic;
  signal core_full: std_logic;
  signal core_dcount: std_logic_vector(data_count_width - 1 downto 0);
begin
  comp0: if ((core_name0 = "fifo_fg92_6a1156e8dc43a711")) generate
    core_instance0: fifo_fg92_6a1156e8dc43a711
      port map (
        clk => clk,
        srst => srst,
        din => din,
        wr_en => wr_en,
        rd_en => rd_en,
        dout => dout,
        full => core_full,
        empty => empty,
        data_count => core_dcount
      );
  end generate;

  modify_count: process(core_full, core_dcount) is
  begin
    if core_full = '1' then
      percent_full <= (others => '1');
    else
      percent_full <= core_dcount(data_count_width-1 downto data_count_width-percent_full_width);
    end if;
  end process modify_count;

  rd_en <= re and en and re_ce;
  wr_en <= we and en and we_ce;
  full <= core_full;
  srst <= rst and ce;
  dcount <= core_dcount;

  terminate_core_ae: if has_ae /= 1 generate
  begin
    ae <= '0';
  end generate terminate_core_ae;
  terminate_core_af: if has_af /= 1 generate
  begin
    af <= '0';
  end generate terminate_core_af;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6dad3a03fc is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6dad3a03fc;


architecture behavior of relational_6dad3a03fc is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_12_17: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 8, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0512fd5e4c is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0512fd5e4c;


architecture behavior of constant_0512fd5e4c is
begin
  op <= "100111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_82fb466a8b is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_82fb466a8b;


architecture behavior of relational_82fb466a8b is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlmult_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    a_width: integer := 4;
    a_bin_pt: integer := 2;
    a_arith: integer := xlSigned;
    b_width: integer := 4;
    b_bin_pt: integer := 1;
    b_arith: integer := xlSigned;
    p_width: integer := 8;
    p_bin_pt: integer := 2;
    p_arith: integer := xlSigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    extra_registers: integer := 0;
    c_a_width: integer := 7;
    c_b_width: integer := 7;
    c_type: integer := 0;
    c_a_type: integer := 0;
    c_b_type: integer := 0;
    c_pipelined: integer := 1;
    c_baat: integer := 4;
    multsign: integer := xlSigned;
    c_output_width: integer := 16
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    core_ce: in std_logic := '0';
    core_clr: in std_logic := '0';
    core_clk: in std_logic := '0';
    rst: in std_logic_vector(rst_width - 1 downto 0);
    en: in std_logic_vector(en_width - 1 downto 0);
    p: out std_logic_vector(p_width - 1 downto 0)
  );
end xlmult_wlan_phy_tx_pmd;
architecture behavior of xlmult_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component mult_11_2_f2bb5a57782af7d9
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of mult_11_2_f2bb5a57782af7d9:
    component is true;
  attribute fpga_dont_touch of mult_11_2_f2bb5a57782af7d9:
    component is "true";
  attribute box_type of mult_11_2_f2bb5a57782af7d9:
    component  is "black_box";
  component mult_11_2_414c0fa5acc33f35
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of mult_11_2_414c0fa5acc33f35:
    component is true;
  attribute fpga_dont_touch of mult_11_2_414c0fa5acc33f35:
    component is "true";
  attribute box_type of mult_11_2_414c0fa5acc33f35:
    component  is "black_box";
  signal tmp_a: std_logic_vector(c_a_width - 1 downto 0);
  signal conv_a: std_logic_vector(c_a_width - 1 downto 0);
  signal tmp_b: std_logic_vector(c_b_width - 1 downto 0);
  signal conv_b: std_logic_vector(c_b_width - 1 downto 0);
  signal tmp_p: std_logic_vector(c_output_width - 1 downto 0);
  signal conv_p: std_logic_vector(p_width - 1 downto 0);
  -- synopsys translate_off
  signal real_a, real_b, real_p: real;
  -- synopsys translate_on
  signal rfd: std_logic;
  signal rdy: std_logic;
  signal nd: std_logic;
  signal internal_ce: std_logic;
  signal internal_clr: std_logic;
  signal internal_core_ce: std_logic;
begin
-- synopsys translate_off
-- synopsys translate_on
  internal_ce <= ce and en(0);
  internal_core_ce <= core_ce and en(0);
  internal_clr <= (clr or rst(0)) and ce;
  nd <= internal_ce;
  input_process:  process (a,b)
  begin
    tmp_a <= zero_ext(a, c_a_width);
    tmp_b <= zero_ext(b, c_b_width);
  end process;
  output_process: process (tmp_p)
  begin
    conv_p <= convert_type(tmp_p, c_output_width, a_bin_pt+b_bin_pt, multsign,
                           p_width, p_bin_pt, p_arith, quantization, overflow);
  end process;
  comp0: if ((core_name0 = "mult_11_2_f2bb5a57782af7d9")) generate
    core_instance0: mult_11_2_f2bb5a57782af7d9
      port map (
        a => tmp_a,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  comp1: if ((core_name0 = "mult_11_2_414c0fa5acc33f35")) generate
    core_instance1: mult_11_2_414c0fa5acc33f35
      port map (
        a => tmp_a,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  latency_gt_0: if (extra_registers > 0) generate
    reg: synth_reg
      generic map (
        width => p_width,
        latency => extra_registers
      )
      port map (
        i => conv_p,
        ce => internal_ce,
        clr => internal_clr,
        clk => clk,
        o => p
      );
  end generate;
  latency_eq_0: if (extra_registers = 0) generate
    p <= conv_p;
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_a54904b290 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((16 - 1) downto 0);
    d1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_a54904b290;


architecture behavior of mux_a54904b290 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((16 - 1) downto 0);
  signal d1_1_27: std_logic_vector((16 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((16 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e25f797841 is
  port (
    in0 : in std_logic_vector((31 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e25f797841;


architecture behavior of concat_e25f797841 is
  signal in0_1_23: unsigned((31 - 1) downto 0);
  signal in1_1_27: boolean;
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= ((in1) = "1");
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & boolean_to_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_bc7a810978 is
  port (
    op : out std_logic_vector((31 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_bc7a810978;


architecture behavior of constant_bc7a810978 is
begin
  op <= "0000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_ddc3ebdd7c is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_ddc3ebdd7c;


architecture behavior of reinterpret_ddc3ebdd7c is
  signal input_port_1_40: unsigned((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_e83dd85005 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_e83dd85005;


architecture behavior of relational_e83dd85005 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1d1da8e0e2 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((3 - 1) downto 0);
    d1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1d1da8e0e2;


architecture behavior of mux_1d1da8e0e2 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((3 - 1) downto 0);
  signal d1_1_27: std_logic_vector((3 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((3 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f9c0f11a18 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((4 - 1) downto 0);
    d1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f9c0f11a18;


architecture behavior of mux_f9c0f11a18 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((4 - 1) downto 0);
  signal d1_1_27: std_logic_vector((4 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((4 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_3e1f051fb7 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_3e1f051fb7;


architecture behavior of logical_3e1f051fb7 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_18f2e784b5 is
  port (
    op : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_18f2e784b5;


architecture behavior of constant_18f2e784b5 is
begin
  op <= "0000001011101001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1e3d9a52c0 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1e3d9a52c0;


architecture behavior of constant_1e3d9a52c0 is
begin
  op <= "00010100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_e55f8c5d80 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((16 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_e55f8c5d80;


architecture behavior of relational_e55f8c5d80 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((16 - 1) downto 0);
  signal cast_22_12: unsigned((16 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_12 <= u2u_cast(a_1_31, 0, 16, 0);
  result_22_3_rel <= cast_22_12 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_60871c3374 is
  port (
    a : in std_logic_vector((5 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_60871c3374;


architecture behavior of relational_60871c3374 is
  signal a_1_31: unsigned((5 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal cast_22_12: unsigned((8 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_22_12 <= u2u_cast(a_1_31, 0, 8, 0);
  result_22_3_rel <= cast_22_12 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_112ed141f4 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_112ed141f4;


architecture behavior of mux_112ed141f4 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((1 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/EDK Processor"

entity edk_processor_entity_de00edcbbe is
  port (
    axi_aresetn: in std_logic; 
    from_register: in std_logic_vector(31 downto 0); 
    plb_ce_1: in std_logic; 
    plb_clk_1: in std_logic; 
    s_axi_araddr: in std_logic_vector(31 downto 0); 
    s_axi_arburst: in std_logic_vector(1 downto 0); 
    s_axi_arcache: in std_logic_vector(3 downto 0); 
    s_axi_arid: in std_logic_vector(7 downto 0); 
    s_axi_arlen: in std_logic_vector(7 downto 0); 
    s_axi_arlock: in std_logic_vector(1 downto 0); 
    s_axi_arprot: in std_logic_vector(2 downto 0); 
    s_axi_arsize: in std_logic_vector(2 downto 0); 
    s_axi_arvalid: in std_logic; 
    s_axi_awaddr: in std_logic_vector(31 downto 0); 
    s_axi_awburst: in std_logic_vector(1 downto 0); 
    s_axi_awcache: in std_logic_vector(3 downto 0); 
    s_axi_awid: in std_logic_vector(7 downto 0); 
    s_axi_awlen: in std_logic_vector(7 downto 0); 
    s_axi_awlock: in std_logic_vector(1 downto 0); 
    s_axi_awprot: in std_logic_vector(2 downto 0); 
    s_axi_awsize: in std_logic_vector(2 downto 0); 
    s_axi_awvalid: in std_logic; 
    s_axi_bready: in std_logic; 
    s_axi_rready: in std_logic; 
    s_axi_wdata: in std_logic_vector(31 downto 0); 
    s_axi_wlast: in std_logic; 
    s_axi_wstrb: in std_logic_vector(3 downto 0); 
    s_axi_wvalid: in std_logic; 
    to_register: in std_logic_vector(31 downto 0); 
    to_register1: in std_logic_vector(31 downto 0); 
    to_register2: in std_logic_vector(31 downto 0); 
    to_register3: in std_logic_vector(31 downto 0); 
    to_register4: in std_logic_vector(31 downto 0); 
    to_register5: in std_logic_vector(31 downto 0); 
    memmap_x0: out std_logic; 
    memmap_x1: out std_logic; 
    memmap_x10: out std_logic; 
    memmap_x11: out std_logic_vector(31 downto 0); 
    memmap_x12: out std_logic; 
    memmap_x13: out std_logic_vector(31 downto 0); 
    memmap_x14: out std_logic; 
    memmap_x15: out std_logic_vector(31 downto 0); 
    memmap_x16: out std_logic; 
    memmap_x17: out std_logic_vector(31 downto 0); 
    memmap_x18: out std_logic; 
    memmap_x19: out std_logic_vector(31 downto 0); 
    memmap_x2: out std_logic_vector(7 downto 0); 
    memmap_x20: out std_logic; 
    memmap_x21: out std_logic_vector(31 downto 0); 
    memmap_x22: out std_logic; 
    memmap_x3: out std_logic_vector(1 downto 0); 
    memmap_x4: out std_logic; 
    memmap_x5: out std_logic_vector(31 downto 0); 
    memmap_x6: out std_logic_vector(7 downto 0); 
    memmap_x7: out std_logic; 
    memmap_x8: out std_logic_vector(1 downto 0); 
    memmap_x9: out std_logic
  );
end edk_processor_entity_de00edcbbe;

architecture structural of edk_processor_entity_de00edcbbe is
  signal axi_aresetn_net_x0: std_logic;
  signal from_register_data_out_net_x0: std_logic_vector(31 downto 0);
  signal memmap_s_axi_arready_net_x0: std_logic;
  signal memmap_s_axi_awready_net_x0: std_logic;
  signal memmap_s_axi_bid_net_x0: std_logic_vector(7 downto 0);
  signal memmap_s_axi_bresp_net_x0: std_logic_vector(1 downto 0);
  signal memmap_s_axi_bvalid_net_x0: std_logic;
  signal memmap_s_axi_rdata_net_x0: std_logic_vector(31 downto 0);
  signal memmap_s_axi_rid_net_x0: std_logic_vector(7 downto 0);
  signal memmap_s_axi_rlast_net_x0: std_logic;
  signal memmap_s_axi_rresp_net_x0: std_logic_vector(1 downto 0);
  signal memmap_s_axi_rvalid_net_x0: std_logic;
  signal memmap_s_axi_wready_net_x0: std_logic;
  signal memmap_sm_config_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_config_en_net_x0: std_logic;
  signal memmap_sm_fft_config_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_fft_config_en_net_x0: std_logic;
  signal memmap_sm_output_scaling_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_output_scaling_en_net_x0: std_logic;
  signal memmap_sm_pkt_buf_sel_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_pkt_buf_sel_en_net_x0: std_logic;
  signal memmap_sm_timing_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_timing_en_net_x0: std_logic;
  signal memmap_sm_tx_start_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_tx_start_en_net_x0: std_logic;
  signal plb_ce_1_sg_x0: std_logic;
  signal plb_clk_1_sg_x0: std_logic;
  signal s_axi_araddr_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_arburst_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_arcache_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_arid_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_arlen_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_arlock_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_arprot_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_arsize_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_arvalid_net_x0: std_logic;
  signal s_axi_awaddr_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_awburst_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_awcache_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_awid_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_awlen_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_awlock_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_awprot_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_awsize_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_awvalid_net_x0: std_logic;
  signal s_axi_bready_net_x0: std_logic;
  signal s_axi_rready_net_x0: std_logic;
  signal s_axi_wdata_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_wlast_net_x0: std_logic;
  signal s_axi_wstrb_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_wvalid_net_x0: std_logic;
  signal to_register1_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register2_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register3_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register4_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register5_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register_dout_net_x0: std_logic_vector(31 downto 0);

begin
  axi_aresetn_net_x0 <= axi_aresetn;
  from_register_data_out_net_x0 <= from_register;
  plb_ce_1_sg_x0 <= plb_ce_1;
  plb_clk_1_sg_x0 <= plb_clk_1;
  s_axi_araddr_net_x0 <= s_axi_araddr;
  s_axi_arburst_net_x0 <= s_axi_arburst;
  s_axi_arcache_net_x0 <= s_axi_arcache;
  s_axi_arid_net_x0 <= s_axi_arid;
  s_axi_arlen_net_x0 <= s_axi_arlen;
  s_axi_arlock_net_x0 <= s_axi_arlock;
  s_axi_arprot_net_x0 <= s_axi_arprot;
  s_axi_arsize_net_x0 <= s_axi_arsize;
  s_axi_arvalid_net_x0 <= s_axi_arvalid;
  s_axi_awaddr_net_x0 <= s_axi_awaddr;
  s_axi_awburst_net_x0 <= s_axi_awburst;
  s_axi_awcache_net_x0 <= s_axi_awcache;
  s_axi_awid_net_x0 <= s_axi_awid;
  s_axi_awlen_net_x0 <= s_axi_awlen;
  s_axi_awlock_net_x0 <= s_axi_awlock;
  s_axi_awprot_net_x0 <= s_axi_awprot;
  s_axi_awsize_net_x0 <= s_axi_awsize;
  s_axi_awvalid_net_x0 <= s_axi_awvalid;
  s_axi_bready_net_x0 <= s_axi_bready;
  s_axi_rready_net_x0 <= s_axi_rready;
  s_axi_wdata_net_x0 <= s_axi_wdata;
  s_axi_wlast_net_x0 <= s_axi_wlast;
  s_axi_wstrb_net_x0 <= s_axi_wstrb;
  s_axi_wvalid_net_x0 <= s_axi_wvalid;
  to_register_dout_net_x0 <= to_register;
  to_register1_dout_net_x0 <= to_register1;
  to_register2_dout_net_x0 <= to_register2;
  to_register3_dout_net_x0 <= to_register3;
  to_register4_dout_net_x0 <= to_register4;
  to_register5_dout_net_x0 <= to_register5;
  memmap_x0 <= memmap_s_axi_arready_net_x0;
  memmap_x1 <= memmap_s_axi_awready_net_x0;
  memmap_x10 <= memmap_s_axi_wready_net_x0;
  memmap_x11 <= memmap_sm_timing_din_net_x0;
  memmap_x12 <= memmap_sm_timing_en_net_x0;
  memmap_x13 <= memmap_sm_config_din_net_x0;
  memmap_x14 <= memmap_sm_config_en_net_x0;
  memmap_x15 <= memmap_sm_pkt_buf_sel_din_net_x0;
  memmap_x16 <= memmap_sm_pkt_buf_sel_en_net_x0;
  memmap_x17 <= memmap_sm_output_scaling_din_net_x0;
  memmap_x18 <= memmap_sm_output_scaling_en_net_x0;
  memmap_x19 <= memmap_sm_tx_start_din_net_x0;
  memmap_x2 <= memmap_s_axi_bid_net_x0;
  memmap_x20 <= memmap_sm_tx_start_en_net_x0;
  memmap_x21 <= memmap_sm_fft_config_din_net_x0;
  memmap_x22 <= memmap_sm_fft_config_en_net_x0;
  memmap_x3 <= memmap_s_axi_bresp_net_x0;
  memmap_x4 <= memmap_s_axi_bvalid_net_x0;
  memmap_x5 <= memmap_s_axi_rdata_net_x0;
  memmap_x6 <= memmap_s_axi_rid_net_x0;
  memmap_x7 <= memmap_s_axi_rlast_net_x0;
  memmap_x8 <= memmap_s_axi_rresp_net_x0;
  memmap_x9 <= memmap_s_axi_rvalid_net_x0;

  memmap: entity work.axi_sgiface
    port map (
      axi_aclk => plb_clk_1_sg_x0,
      axi_aresetn => axi_aresetn_net_x0,
      axi_ce => plb_ce_1_sg_x0,
      s_axi_araddr => s_axi_araddr_net_x0,
      s_axi_arburst => s_axi_arburst_net_x0,
      s_axi_arcache => s_axi_arcache_net_x0,
      s_axi_arid => s_axi_arid_net_x0,
      s_axi_arlen => s_axi_arlen_net_x0,
      s_axi_arlock => s_axi_arlock_net_x0,
      s_axi_arprot => s_axi_arprot_net_x0,
      s_axi_arsize => s_axi_arsize_net_x0,
      s_axi_arvalid => s_axi_arvalid_net_x0,
      s_axi_awaddr => s_axi_awaddr_net_x0,
      s_axi_awburst => s_axi_awburst_net_x0,
      s_axi_awcache => s_axi_awcache_net_x0,
      s_axi_awid => s_axi_awid_net_x0,
      s_axi_awlen => s_axi_awlen_net_x0,
      s_axi_awlock => s_axi_awlock_net_x0,
      s_axi_awprot => s_axi_awprot_net_x0,
      s_axi_awsize => s_axi_awsize_net_x0,
      s_axi_awvalid => s_axi_awvalid_net_x0,
      s_axi_bready => s_axi_bready_net_x0,
      s_axi_rready => s_axi_rready_net_x0,
      s_axi_wdata => s_axi_wdata_net_x0,
      s_axi_wlast => s_axi_wlast_net_x0,
      s_axi_wstrb => s_axi_wstrb_net_x0,
      s_axi_wvalid => s_axi_wvalid_net_x0,
      sm_config_dout => to_register1_dout_net_x0,
      sm_fft_config_dout => to_register5_dout_net_x0,
      sm_output_scaling_dout => to_register3_dout_net_x0,
      sm_pkt_buf_sel_dout => to_register2_dout_net_x0,
      sm_status_dout => from_register_data_out_net_x0,
      sm_timing_dout => to_register_dout_net_x0,
      sm_tx_start_dout => to_register4_dout_net_x0,
      s_axi_arready => memmap_s_axi_arready_net_x0,
      s_axi_awready => memmap_s_axi_awready_net_x0,
      s_axi_bid => memmap_s_axi_bid_net_x0,
      s_axi_bresp => memmap_s_axi_bresp_net_x0,
      s_axi_bvalid => memmap_s_axi_bvalid_net_x0,
      s_axi_rdata => memmap_s_axi_rdata_net_x0,
      s_axi_rid => memmap_s_axi_rid_net_x0,
      s_axi_rlast => memmap_s_axi_rlast_net_x0,
      s_axi_rresp => memmap_s_axi_rresp_net_x0,
      s_axi_rvalid => memmap_s_axi_rvalid_net_x0,
      s_axi_wready => memmap_s_axi_wready_net_x0,
      sm_config_din => memmap_sm_config_din_net_x0,
      sm_config_en => memmap_sm_config_en_net_x0,
      sm_fft_config_din => memmap_sm_fft_config_din_net_x0,
      sm_fft_config_en => memmap_sm_fft_config_en_net_x0,
      sm_output_scaling_din => memmap_sm_output_scaling_din_net_x0,
      sm_output_scaling_en => memmap_sm_output_scaling_en_net_x0,
      sm_pkt_buf_sel_din => memmap_sm_pkt_buf_sel_din_net_x0,
      sm_pkt_buf_sel_en => memmap_sm_pkt_buf_sel_en_net_x0,
      sm_timing_din => memmap_sm_timing_din_net_x0,
      sm_timing_en => memmap_sm_timing_en_net_x0,
      sm_tx_start_din => memmap_sm_tx_start_din_net_x0,
      sm_tx_start_en => memmap_sm_tx_start_en_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/HT Preamble Gen/S-R Latch1"

entity s_r_latch1_entity_18268c34fe is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    r: in std_logic; 
    s: in std_logic; 
    q: out std_logic
  );
end s_r_latch1_entity_18268c34fe;

architecture structural of s_r_latch1_entity_18268c34fe is
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant1_op_net: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;

begin
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  logical2_y_net_x0 <= r;
  logical3_y_net_x0 <= s;
  q <= register2_q_net_x0;

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => logical2_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => logical3_y_net_x0,
      en => "1",
      dout(0) => convert2_dout_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => constant1_op_net,
      en(0) => convert2_dout_net,
      rst(0) => convert1_dout_net,
      q(0) => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/HT Preamble Gen"

entity ht_preamble_gen_entity_624eef30fb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    iq_fifo_tready: in std_logic; 
    start: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    tx_reset: in std_logic; 
    delay1_x0: out std_logic; 
    delay2_x0: out std_logic; 
    ht_training_q_x0: out std_logic_vector(15 downto 0); 
    iq_stream: out std_logic_vector(15 downto 0); 
    sym_cfg_x0: out std_logic_vector(17 downto 0)
  );
end ht_preamble_gen_entity_624eef30fb;

architecture structural of ht_preamble_gen_entity_624eef30fb is
  signal axi_fifo_s_axis_tready_net_x0: std_logic;
  signal ce_1_sg_x1: std_logic;
  signal clk_1_sg_x1: std_logic;
  signal concat_y_net: std_logic_vector(6 downto 0);
  signal concat_y_net_x1: std_logic_vector(17 downto 0);
  signal constant9_op_net: std_logic_vector(5 downto 0);
  signal counter1_op_net: std_logic_vector(5 downto 0);
  signal delay3_q_net: std_logic;
  signal delay_q_net_x0: std_logic_vector(17 downto 0);
  signal i_x0: std_logic_vector(15 downto 0);
  signal inverter1_op_net: std_logic;
  signal iq_tlast_x0: std_logic;
  signal iq_tvalid_x0: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical4_y_net: std_logic;
  signal logical4_y_net_x1: std_logic;
  signal logical_y_net_x0: std_logic;
  signal mcode_load_htltf_net: std_logic;
  signal mcode_load_htstf_net: std_logic;
  signal q_x0: std_logic_vector(15 downto 0);
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;

begin
  ce_1_sg_x1 <= ce_1;
  clk_1_sg_x1 <= clk_1;
  axi_fifo_s_axis_tready_net_x0 <= iq_fifo_tready;
  logical4_y_net_x1 <= start;
  concat_y_net_x1 <= sym_cfg;
  logical_y_net_x0 <= tx_reset;
  delay1_x0 <= iq_tvalid_x0;
  delay2_x0 <= iq_tlast_x0;
  ht_training_q_x0 <= q_x0;
  iq_stream <= i_x0;
  sym_cfg_x0 <= delay_q_net_x0;

  concat: entity work.concat_0d20f96564
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay3_q_net,
      in1 => counter1_op_net,
      y => concat_y_net
    );

  constant9: entity work.constant_c462ec0feb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant9_op_net
    );

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_f068fb73312ae1e5",
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      clr => '0',
      en(0) => logical4_y_net,
      rst(0) => inverter1_op_net,
      op => counter1_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      d => concat_y_net_x1,
      en => '1',
      rst => '1',
      q => delay_q_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => iq_tvalid_x0
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      d(0) => relational2_op_net,
      en => '1',
      rst => '1',
      q(0) => iq_tlast_x0
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      d(0) => mcode_load_htltf_net,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net
    );

  ht_training_i: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 7,
      c_address_width => 7,
      c_width => 16,
      core_name0 => "dmg_72_48a0132db6517610",
      latency => 1
    )
    port map (
      addr => concat_y_net,
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      en => "1",
      data => i_x0
    );

  ht_training_q: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 7,
      c_address_width => 7,
      c_width => 16,
      core_name0 => "dmg_72_2be916f69ff4e5b8",
      latency => 1
    )
    port map (
      addr => concat_y_net,
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      en => "1",
      data => q_x0
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => mcode_load_htltf_net,
      d1(0) => mcode_load_htstf_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x0,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net,
      d1(0) => logical4_y_net_x1,
      y(0) => logical3_y_net_x0
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => axi_fifo_s_axis_tready_net_x0,
      y(0) => logical4_y_net
    );

  mcode: entity work.mcode_block_00412594a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      sym_cfg => concat_y_net_x1,
      load_htltf(0) => mcode_load_htltf_net,
      load_htstf(0) => mcode_load_htstf_net
    );

  relational2: entity work.relational_15ce3046b2
    port map (
      a => counter1_op_net,
      b => constant9_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  s_r_latch1_18268c34fe: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x1,
      clk_1 => clk_1_sg_x1,
      r => logical2_y_net_x0,
      s => logical3_y_net_x0,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/Buffer and Cyclic Prefix/Control"

entity control_entity_3a56a32023 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    regtx_cp_len: in std_logic_vector(7 downto 0); 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    tlast: in std_logic; 
    rd_addr: out std_logic_vector(7 downto 0); 
    valid: out std_logic
  );
end control_entity_3a56a32023;

architecture structural of control_entity_3a56a32023 is
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal ce_1_sg_x3: std_logic;
  signal clk_1_sg_x3: std_logic;
  signal counter_op_net_x0: std_logic_vector(7 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x1: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register8_q_net_x0: std_logic_vector(7 downto 0);
  signal register9_q_net_x0: std_logic_vector(7 downto 0);
  signal relational3_op_net_x0: std_logic;

begin
  ce_1_sg_x3 <= ce_1;
  clk_1_sg_x3 <= clk_1;
  register9_q_net_x0 <= regtx_cp_len;
  register8_q_net_x0 <= regtx_num_sc;
  fast_fourier_transform_8_0_m_axis_data_tlast_net_x1 <= tlast;
  rd_addr <= counter_op_net_x0;
  valid <= logical2_y_net_x0;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 8,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 9,
      core_name0 => "addsb_11_0_60fd3b5996582b7a",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 9,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => register8_q_net_x0,
      b => register9_q_net_x0,
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_86806e294f737f4c",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      clr => '0',
      en(0) => register2_q_net_x0,
      rst(0) => inverter1_op_net,
      op => counter_op_net_x0
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      clr => '0',
      ip(0) => relational3_op_net_x0,
      op(0) => inverter2_op_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => inverter2_op_net,
      y(0) => logical2_y_net_x0
    );

  relational3: entity work.relational_305a9068e6
    port map (
      a => counter_op_net_x0,
      b => addsub_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net_x0
    );

  s_r_latch1_c008c4d1e2: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x3,
      clk_1 => clk_1_sg_x3,
      r => relational3_op_net_x0,
      s => fast_fourier_transform_8_0_m_axis_data_tlast_net_x1,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/Buffer and Cyclic Prefix/I/Q Concat"

entity q_concat_entity_4cbb243c07 is
  port (
    i: in std_logic_vector(15 downto 0); 
    q: in std_logic_vector(15 downto 0); 
    iq: out std_logic_vector(31 downto 0)
  );
end q_concat_entity_4cbb243c07;

architecture structural of q_concat_entity_4cbb243c07 is
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0 <= i;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0 <= q;
  iq <= concat_y_net_x0;

  concat: entity work.concat_a369e00c6b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net_x0
    );

  reinterpret: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/Buffer and Cyclic Prefix/I/Q Slice"

entity q_slice_entity_6da961fd0c is
  port (
    iq: in std_logic_vector(31 downto 0); 
    i: out std_logic_vector(15 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end q_slice_entity_6da961fd0c;

architecture structural of q_slice_entity_6da961fd0c is
  signal dual_port_ram_doutb_net_x0: std_logic_vector(31 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(15 downto 0);
  signal slice1_y_net: std_logic_vector(15 downto 0);
  signal slice_y_net: std_logic_vector(15 downto 0);

begin
  dual_port_ram_doutb_net_x0 <= iq;
  i <= reinterpret2_output_port_net_x0;
  q <= reinterpret3_output_port_net_x0;

  reinterpret2: entity work.reinterpret_151459306d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_151459306d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 31,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => dual_port_ram_doutb_net_x0,
      y => slice_y_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 15,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => dual_port_ram_doutb_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/Buffer and Cyclic Prefix"

entity buffer_and_cyclic_prefix_entity_435e2544cb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    q: in std_logic_vector(15 downto 0); 
    regtx_cp_len: in std_logic_vector(7 downto 0); 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    tlast: in std_logic; 
    tvalid: in std_logic; 
    xkindex: in std_logic_vector(5 downto 0); 
    i_x0: out std_logic_vector(15 downto 0); 
    q_x0: out std_logic_vector(15 downto 0); 
    valid: out std_logic
  );
end buffer_and_cyclic_prefix_entity_435e2544cb;

architecture structural of buffer_and_cyclic_prefix_entity_435e2544cb is
  signal addsub1_s_net: std_logic_vector(5 downto 0);
  signal addsub2_s_net: std_logic_vector(8 downto 0);
  signal ce_1_sg_x4: std_logic;
  signal clk_1_sg_x4: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant1_op_net: std_logic_vector(31 downto 0);
  signal constant2_op_net: std_logic;
  signal counter_op_net_x0: std_logic_vector(7 downto 0);
  signal delay3_q_net_x0: std_logic;
  signal dual_port_ram_doutb_net_x0: std_logic_vector(31 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x2: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x0: std_logic_vector(5 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal register8_q_net_x1: std_logic_vector(7 downto 0);
  signal register9_q_net_x1: std_logic_vector(7 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x4 <= ce_1;
  clk_1_sg_x4 <= clk_1;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1 <= i;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1 <= q;
  register9_q_net_x1 <= regtx_cp_len;
  register8_q_net_x1 <= regtx_num_sc;
  fast_fourier_transform_8_0_m_axis_data_tlast_net_x2 <= tlast;
  fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0 <= tvalid;
  fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x0 <= xkindex;
  i_x0 <= reinterpret2_output_port_net_x1;
  q_x0 <= reinterpret3_output_port_net_x1;
  valid <= delay3_q_net_x0;

  addsub1: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 0,
      a_width => 9,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 8,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 10,
      core_name0 => "addsb_11_0_d5bf78f2384e976c",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 10,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 6
    )
    port map (
      a => addsub2_s_net,
      b => counter_op_net_x0,
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      en => "1",
      s => addsub1_s_net
    );

  addsub2: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 8,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 9,
      core_name0 => "addsb_11_0_8942e2ad5d8d4897",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 9,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => register8_q_net_x1,
      b => register9_q_net_x1,
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      en => "1",
      s => addsub2_s_net
    );

  constant1: entity work.constant_37567836aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  control_3a56a32023: entity work.control_entity_3a56a32023
    port map (
      ce_1 => ce_1_sg_x4,
      clk_1 => clk_1_sg_x4,
      regtx_cp_len => register9_q_net_x1,
      regtx_num_sc => register8_q_net_x1,
      tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x2,
      rd_addr => counter_op_net_x0,
      valid => logical2_y_net_x0
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      d(0) => logical2_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x0
    );

  dual_port_ram: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 6,
      c_address_width_b => 6,
      c_width_a => 32,
      c_width_b => 32,
      core_name0 => "bmg_72_e4abe4c74ea5aa02",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x4,
      a_clk => clk_1_sg_x4,
      addra => fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x0,
      addrb => addsub1_s_net,
      b_ce => ce_1_sg_x4,
      b_clk => clk_1_sg_x4,
      dina => concat_y_net_x0,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0,
      web(0) => constant2_op_net,
      doutb => dual_port_ram_doutb_net_x0
    );

  q_concat_4cbb243c07: entity work.q_concat_entity_4cbb243c07
    port map (
      i => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1,
      q => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1,
      iq => concat_y_net_x0
    );

  q_slice_6da961fd0c: entity work.q_slice_entity_6da961fd0c
    port map (
      iq => dual_port_ram_doutb_net_x0,
      i => reinterpret2_output_port_net_x1,
      q => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/FFT Core"

entity fft_core_entity_2954b1083d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    iq_in_valid: in std_logic; 
    iq_tlast: in std_logic; 
    q: in std_logic_vector(15 downto 0); 
    regtx_fft_scaling: in std_logic_vector(5 downto 0); 
    tx_reset: in std_logic; 
    data_in_tready: out std_logic; 
    data_out_tlast: out std_logic; 
    data_out_tvalid: out std_logic; 
    data_xk_index: out std_logic_vector(5 downto 0); 
    i_out: out std_logic_vector(15 downto 0); 
    q_out: out std_logic_vector(15 downto 0)
  );
end fft_core_entity_2954b1083d;

architecture structural of fft_core_entity_2954b1083d is
  signal axi_fifo_m_axis_tvalid_net_x0: std_logic;
  signal ce_1_sg_x5: std_logic;
  signal clk_1_sg_x5: std_logic;
  signal constant1_op_net: std_logic;
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant4_op_net: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x3: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1: std_logic_vector(5 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x0: std_logic;
  signal inverter_op_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x1: std_logic;
  signal register10_q_net_x0: std_logic_vector(5 downto 0);
  signal register_q_net: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x5 <= ce_1;
  clk_1_sg_x5 <= clk_1;
  reinterpret2_output_port_net_x0 <= i;
  axi_fifo_m_axis_tvalid_net_x0 <= iq_in_valid;
  logical2_y_net_x0 <= iq_tlast;
  reinterpret3_output_port_net_x0 <= q;
  register10_q_net_x0 <= regtx_fft_scaling;
  logical_y_net_x1 <= tx_reset;
  data_in_tready <= fast_fourier_transform_8_0_s_axis_data_tready_net_x0;
  data_out_tlast <= fast_fourier_transform_8_0_m_axis_data_tlast_net_x3;
  data_out_tvalid <= fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1;
  data_xk_index <= fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1;
  i_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2;
  q_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant2: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant4: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant4_op_net
    );

  fast_fourier_transform_8_0: entity work.xlfast_fourier_transform_886093b6a909385035fdd94c865209c9
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      m_axis_data_tready => constant3_op_net,
      m_axis_status_tready => constant2_op_net,
      rst => register_q_net,
      s_axis_config_tdata_fwd_inv(0) => constant1_op_net,
      s_axis_config_tdata_scale_sch => register10_q_net_x0,
      s_axis_config_tvalid => constant4_op_net,
      s_axis_data_tdata_xn_im => reinterpret3_output_port_net_x0,
      s_axis_data_tdata_xn_re => reinterpret2_output_port_net_x0,
      s_axis_data_tlast => logical2_y_net_x0,
      s_axis_data_tvalid => axi_fifo_m_axis_tvalid_net_x0,
      m_axis_data_tdata_xk_im => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2,
      m_axis_data_tdata_xk_re => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2,
      m_axis_data_tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x3,
      m_axis_data_tuser_xk_index => fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1,
      m_axis_data_tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1,
      s_axis_data_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x0
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      clr => '0',
      ip(0) => logical_y_net_x1,
      op(0) => inverter_op_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      d(0) => inverter_op_net,
      en => "1",
      rst => "0",
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix/FIFO"

entity fifo_entity_c7741c9113 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_tready: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    iq_tlast: in std_logic; 
    iq_tvalid: in std_logic; 
    q: in std_logic_vector(15 downto 0); 
    sym_cfg: in std_logic_vector(17 downto 0); 
    tx_reset: in std_logic; 
    fifo_tready: out std_logic; 
    i_x0: out std_logic_vector(15 downto 0); 
    iq_tlast_x0: out std_logic; 
    iq_tvalid_x0: out std_logic; 
    q_x0: out std_logic_vector(15 downto 0)
  );
end fifo_entity_c7741c9113;

architecture structural of fifo_entity_c7741c9113 is
  signal axi_fifo_m_axis_tdata_net_x0: std_logic_vector(31 downto 0);
  signal axi_fifo_m_axis_tlast_net: std_logic;
  signal axi_fifo_m_axis_tvalid_net_x1: std_logic;
  signal axi_fifo_s_axis_tready_net_x1: std_logic;
  signal ce_1_sg_x6: std_logic;
  signal clk_1_sg_x6: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert1_dout_net_x0: std_logic_vector(15 downto 0);
  signal convert_dout_net_x0: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x1: std_logic;
  signal inverter_op_net: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(15 downto 0);
  signal mux2_y_net_x0: std_logic;
  signal mux3_y_net_x0: std_logic;
  signal mux4_y_net_x0: std_logic_vector(17 downto 0);
  signal mux6_y_net_x0: std_logic_vector(15 downto 0);
  signal register_q_net: std_logic;
  signal reinterpret2_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x6 <= ce_1;
  clk_1_sg_x6 <= clk_1;
  fast_fourier_transform_8_0_s_axis_data_tready_net_x1 <= fft_tready;
  mux6_y_net_x0 <= i;
  mux3_y_net_x0 <= iq_tlast;
  mux2_y_net_x0 <= iq_tvalid;
  mux1_y_net_x0 <= q;
  mux4_y_net_x0 <= sym_cfg;
  logical_y_net_x2 <= tx_reset;
  fifo_tready <= axi_fifo_s_axis_tready_net_x1;
  i_x0 <= reinterpret2_output_port_net_x2;
  iq_tlast_x0 <= logical2_y_net_x1;
  iq_tvalid_x0 <= axi_fifo_m_axis_tvalid_net_x1;
  q_x0 <= reinterpret3_output_port_net_x2;

  axi_fifo: entity work.xlaxififogen_wlan_phy_tx_pmd
    generic map (
      core_name0 => "axififo_fg92_83e0abc99b742965",
      depth_bits => 8,
      has_aresetn => 1,
      tdata_width => 32,
      tuser_width => 18
    )
    port map (
      aresetn => register_q_net,
      ce => ce_1_sg_x6,
      m_axis_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x1,
      s_aclk => clk_1_sg_x6,
      s_axis_tdata => concat_y_net_x0,
      s_axis_tlast => mux3_y_net_x0,
      s_axis_tuser => mux4_y_net_x0,
      s_axis_tvalid => mux2_y_net_x0,
      m_axis_tdata => axi_fifo_m_axis_tdata_net_x0,
      m_axis_tlast => axi_fifo_m_axis_tlast_net,
      m_axis_tvalid => axi_fifo_m_axis_tvalid_net_x1,
      s_axis_tready => axi_fifo_s_axis_tready_net_x1
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      din => mux6_y_net_x0,
      en => "1",
      dout => convert_dout_net_x0
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      din => mux1_y_net_x0,
      en => "1",
      dout => convert1_dout_net_x0
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      ip(0) => logical_y_net_x2,
      op(0) => inverter_op_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => axi_fifo_m_axis_tvalid_net_x1,
      d1(0) => axi_fifo_m_axis_tlast_net,
      y(0) => logical2_y_net_x1
    );

  q_concat_d6adc1378a: entity work.q_concat_entity_4cbb243c07
    port map (
      i => convert_dout_net_x0,
      q => convert1_dout_net_x0,
      iq => concat_y_net_x0
    );

  q_slice_2f21a0a3a6: entity work.q_slice_entity_6da961fd0c
    port map (
      iq => axi_fifo_m_axis_tdata_net_x0,
      i => reinterpret2_output_port_net_x2,
      q => reinterpret3_output_port_net_x2
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      d(0) => inverter_op_net,
      en => "1",
      rst => "0",
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/IFFT and Cyclic Prefix"

entity ifft_and_cyclic_prefix_entity_d9041c6806 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    iq_tlast: in std_logic; 
    iq_valid: in std_logic; 
    logical: in std_logic; 
    q: in std_logic_vector(15 downto 0); 
    register10: in std_logic_vector(5 downto 0); 
    register8: in std_logic_vector(7 downto 0); 
    register9: in std_logic_vector(7 downto 0); 
    sym_cfg: in std_logic_vector(17 downto 0); 
    fifo_tready: out std_logic; 
    i_x0: out std_logic_vector(15 downto 0); 
    iq_valid_x0: out std_logic; 
    q_x0: out std_logic_vector(15 downto 0)
  );
end ifft_and_cyclic_prefix_entity_d9041c6806;

architecture structural of ifft_and_cyclic_prefix_entity_d9041c6806 is
  signal axi_fifo_m_axis_tvalid_net_x1: std_logic;
  signal axi_fifo_s_axis_tready_net_x2: std_logic;
  signal ce_1_sg_x7: std_logic;
  signal clk_1_sg_x7: std_logic;
  signal delay3_q_net_x1: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x3: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1: std_logic_vector(5 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x1: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net_x3: std_logic;
  signal mux1_y_net_x1: std_logic_vector(15 downto 0);
  signal mux2_y_net_x1: std_logic;
  signal mux3_y_net_x1: std_logic;
  signal mux4_y_net_x1: std_logic_vector(17 downto 0);
  signal mux6_y_net_x1: std_logic_vector(15 downto 0);
  signal register10_q_net_x1: std_logic_vector(5 downto 0);
  signal register8_q_net_x2: std_logic_vector(7 downto 0);
  signal register9_q_net_x2: std_logic_vector(7 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x3: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x7 <= ce_1;
  clk_1_sg_x7 <= clk_1;
  mux6_y_net_x1 <= i;
  mux3_y_net_x1 <= iq_tlast;
  mux2_y_net_x1 <= iq_valid;
  logical_y_net_x3 <= logical;
  mux1_y_net_x1 <= q;
  register10_q_net_x1 <= register10;
  register8_q_net_x2 <= register8;
  register9_q_net_x2 <= register9;
  mux4_y_net_x1 <= sym_cfg;
  fifo_tready <= axi_fifo_s_axis_tready_net_x2;
  i_x0 <= reinterpret2_output_port_net_x3;
  iq_valid_x0 <= delay3_q_net_x1;
  q_x0 <= reinterpret3_output_port_net_x3;

  buffer_and_cyclic_prefix_435e2544cb: entity work.buffer_and_cyclic_prefix_entity_435e2544cb
    port map (
      ce_1 => ce_1_sg_x7,
      clk_1 => clk_1_sg_x7,
      i => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2,
      q => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2,
      regtx_cp_len => register9_q_net_x2,
      regtx_num_sc => register8_q_net_x2,
      tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x3,
      tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1,
      xkindex => fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1,
      i_x0 => reinterpret2_output_port_net_x3,
      q_x0 => reinterpret3_output_port_net_x3,
      valid => delay3_q_net_x1
    );

  fft_core_2954b1083d: entity work.fft_core_entity_2954b1083d
    port map (
      ce_1 => ce_1_sg_x7,
      clk_1 => clk_1_sg_x7,
      i => reinterpret2_output_port_net_x2,
      iq_in_valid => axi_fifo_m_axis_tvalid_net_x1,
      iq_tlast => logical2_y_net_x1,
      q => reinterpret3_output_port_net_x2,
      regtx_fft_scaling => register10_q_net_x1,
      tx_reset => logical_y_net_x3,
      data_in_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x1,
      data_out_tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x3,
      data_out_tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1,
      data_xk_index => fast_fourier_transform_8_0_m_axis_data_tuser_xk_index_net_x1,
      i_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2,
      q_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2
    );

  fifo_c7741c9113: entity work.fifo_entity_c7741c9113
    port map (
      ce_1 => ce_1_sg_x7,
      clk_1 => clk_1_sg_x7,
      fft_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x1,
      i => mux6_y_net_x1,
      iq_tlast => mux3_y_net_x1,
      iq_tvalid => mux2_y_net_x1,
      q => mux1_y_net_x1,
      sym_cfg => mux4_y_net_x1,
      tx_reset => logical_y_net_x3,
      fifo_tready => axi_fifo_s_axis_tready_net_x2,
      i_x0 => reinterpret2_output_port_net_x2,
      iq_tlast_x0 => logical2_y_net_x1,
      iq_tvalid_x0 => axi_fifo_m_axis_tvalid_net_x1,
      q_x0 => reinterpret3_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Mux"

entity mux_entity_e0e38b1125 is
  port (
    delay: in std_logic; 
    delay1: in std_logic; 
    ht_preamble_gen: in std_logic; 
    ht_preamble_gen_x0: in std_logic; 
    ht_preamble_gen_x1: in std_logic_vector(15 downto 0); 
    mux4_x0: in std_logic_vector(11 downto 0); 
    preamble_iq: in std_logic_vector(15 downto 0); 
    preamble_sym_cfg: in std_logic_vector(17 downto 0); 
    psdu_iq: in std_logic_vector(11 downto 0); 
    psdu_sym_cfg: in std_logic_vector(17 downto 0); 
    i: out std_logic_vector(15 downto 0); 
    iq_tlast: out std_logic; 
    iq_tvalid: out std_logic; 
    q: out std_logic_vector(15 downto 0); 
    sym_cfg: out std_logic_vector(17 downto 0)
  );
end mux_entity_e0e38b1125;

architecture structural of mux_entity_e0e38b1125 is
  signal delay1_q_net_x0: std_logic;
  signal delay_q_net_x2: std_logic_vector(17 downto 0);
  signal delay_q_net_x3: std_logic;
  signal delay_q_net_x4: std_logic_vector(17 downto 0);
  signal i_x1: std_logic_vector(15 downto 0);
  signal iq_tlast_x1: std_logic;
  signal iq_tvalid_x1: std_logic;
  signal mux1_y_net_x2: std_logic_vector(15 downto 0);
  signal mux2_y_net_x2: std_logic;
  signal mux3_y_net_x0: std_logic_vector(11 downto 0);
  signal mux3_y_net_x2: std_logic;
  signal mux4_y_net_x0: std_logic_vector(11 downto 0);
  signal mux4_y_net_x2: std_logic_vector(17 downto 0);
  signal mux6_y_net_x2: std_logic_vector(15 downto 0);
  signal q_x1: std_logic_vector(15 downto 0);

begin
  delay_q_net_x3 <= delay;
  delay1_q_net_x0 <= delay1;
  iq_tvalid_x1 <= ht_preamble_gen;
  iq_tlast_x1 <= ht_preamble_gen_x0;
  q_x1 <= ht_preamble_gen_x1;
  mux4_y_net_x0 <= mux4_x0;
  i_x1 <= preamble_iq;
  delay_q_net_x2 <= preamble_sym_cfg;
  mux3_y_net_x0 <= psdu_iq;
  delay_q_net_x4 <= psdu_sym_cfg;
  i <= mux6_y_net_x2;
  iq_tlast <= mux3_y_net_x2;
  iq_tvalid <= mux2_y_net_x2;
  q <= mux1_y_net_x2;
  sym_cfg <= mux4_y_net_x2;

  mux1: entity work.mux_35690eb8ec
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => q_x1,
      d1 => mux4_y_net_x0,
      sel(0) => delay_q_net_x3,
      y => mux1_y_net_x2
    );

  mux2: entity work.mux_d99e59b6d4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => iq_tvalid_x1,
      d1(0) => delay_q_net_x3,
      sel(0) => delay_q_net_x3,
      y(0) => mux2_y_net_x2
    );

  mux3: entity work.mux_d99e59b6d4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => iq_tlast_x1,
      d1(0) => delay1_q_net_x0,
      sel(0) => delay_q_net_x3,
      y(0) => mux3_y_net_x2
    );

  mux4: entity work.mux_42c705c90b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => delay_q_net_x2,
      d1 => delay_q_net_x4,
      sel(0) => delay_q_net_x3,
      y => mux4_y_net_x2
    );

  mux6: entity work.mux_35690eb8ec
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => i_x1,
      d1 => mux3_y_net_x0,
      sel(0) => delay_q_net_x3,
      y => mux6_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/OFDM Symbol Ctrl/Posedge1"

entity posedge1_entity_78541e5bea is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end posedge1_entity_78541e5bea;

architecture structural of posedge1_entity_78541e5bea is
  signal ce_1_sg_x8: std_logic;
  signal clk_1_sg_x8: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal register3_q_net_x0: std_logic;

begin
  ce_1_sg_x8 <= ce_1;
  clk_1_sg_x8 <= clk_1;
  register3_q_net_x0 <= d;
  q <= logical1_y_net_x0;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x8,
      clk => clk_1_sg_x8,
      d(0) => register3_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x8,
      clk => clk_1_sg_x8,
      clr => '0',
      ip(0) => delay_q_net,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => register3_q_net_x0,
      y(0) => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/OFDM Symbol Ctrl/Sym Config Encode"

entity sym_config_encode_entity_43a940459d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ofdm_sym_ind: in std_logic_vector(9 downto 0); 
    tx_phy_mode_11ag: in std_logic; 
    tx_phy_mode_11n: in std_logic; 
    tx_phy_mode_11n_ac: in std_logic; 
    sym_cfg: out std_logic_vector(17 downto 0)
  );
end sym_config_encode_entity_43a940459d;

architecture structural of sym_config_encode_entity_43a940459d is
  signal addsub_s_net: std_logic_vector(1 downto 0);
  signal ce_1_sg_x14: std_logic;
  signal clk_1_sg_x14: std_logic;
  signal concat_y_net_x2: std_logic_vector(17 downto 0);
  signal constant10_op_net: std_logic_vector(2 downto 0);
  signal constant11_op_net: std_logic;
  signal constant12_op_net: std_logic_vector(1 downto 0);
  signal constant13_op_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(4 downto 0);
  signal constant2_op_net: std_logic_vector(4 downto 0);
  signal constant3_op_net: std_logic;
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal constant5_op_net: std_logic;
  signal constant6_op_net: std_logic_vector(2 downto 0);
  signal constant7_op_net: std_logic;
  signal constant8_op_net: std_logic_vector(1 downto 0);
  signal constant9_op_net: std_logic_vector(1 downto 0);
  signal logical10_y_net: std_logic;
  signal logical11_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical4_y_net: std_logic;
  signal logical5_y_net: std_logic;
  signal logical6_y_net: std_logic;
  signal logical7_y_net: std_logic;
  signal logical8_y_net: std_logic;
  signal logical9_y_net: std_logic;
  signal mux_y_net: std_logic_vector(1 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational4_op_net: std_logic;
  signal relational5_op_net: std_logic;
  signal relational6_op_net: std_logic;
  signal relational7_op_net: std_logic;
  signal relational_op_net: std_logic;
  signal slice1_y_net_x0: std_logic;
  signal slice_y_net_x0: std_logic;
  signal sym_counter_op_net_x0: std_logic_vector(9 downto 0);
  signal x2lsb_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x14 <= ce_1;
  clk_1_sg_x14 <= clk_1;
  sym_counter_op_net_x0 <= ofdm_sym_ind;
  slice_y_net_x0 <= tx_phy_mode_11ag;
  slice1_y_net_x0 <= tx_phy_mode_11n;
  logical3_y_net_x1 <= tx_phy_mode_11n_ac;
  sym_cfg <= concat_y_net_x2;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_5c670787eb4ba225",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => x2lsb_y_net,
      b => constant13_op_net,
      ce => ce_1_sg_x14,
      clk => clk_1_sg_x14,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  concat: entity work.concat_91ce9c6dac
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant2_op_net,
      in1 => constant1_op_net,
      in2(0) => constant11_op_net,
      in3 => mux_y_net,
      in4(0) => logical5_y_net,
      in5(0) => logical11_y_net,
      in6(0) => logical10_y_net,
      in7(0) => logical8_y_net,
      in8(0) => logical3_y_net,
      y => concat_y_net_x2
    );

  constant1: entity work.constant_ef0e2e5fc6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant10: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant10_op_net
    );

  constant11: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant11_op_net
    );

  constant12: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant12_op_net
    );

  constant13: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant13_op_net
    );

  constant2: entity work.constant_fe72737ca0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant4: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant5_op_net
    );

  constant6: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  constant7: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant7_op_net
    );

  constant8: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net
    );

  constant9: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant9_op_net
    );

  logical10: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational6_op_net,
      d1(0) => slice1_y_net_x0,
      y(0) => logical10_y_net
    );

  logical11: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational7_op_net,
      d1(0) => slice1_y_net_x0,
      y(0) => logical11_y_net
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational_op_net,
      d1(0) => logical4_y_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net,
      d1(0) => logical3_y_net_x1,
      y(0) => logical4_y_net
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical7_y_net,
      d1(0) => logical6_y_net,
      y(0) => logical5_y_net
    );

  logical6: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => slice1_y_net_x0,
      y(0) => logical6_y_net
    );

  logical7: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational2_op_net,
      d1(0) => slice_y_net_x0,
      y(0) => logical7_y_net
    );

  logical8: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical9_y_net,
      d1(0) => slice1_y_net_x0,
      y(0) => logical8_y_net
    );

  logical9: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational4_op_net,
      d1(0) => relational5_op_net,
      y(0) => logical9_y_net
    );

  mux: entity work.mux_2a63ac73aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant12_op_net,
      d1 => addsub_s_net,
      sel(0) => logical6_y_net,
      y => mux_y_net
    );

  relational: entity work.relational_1d0997f32b
    port map (
      a => sym_counter_op_net_x0,
      b(0) => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_0f9b7ba263
    port map (
      a => sym_counter_op_net_x0,
      b => constant4_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_3c449faea2
    port map (
      a => sym_counter_op_net_x0,
      b(0) => constant5_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_7907e32f0f
    port map (
      a => sym_counter_op_net_x0,
      b => constant6_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  relational4: entity work.relational_1d0997f32b
    port map (
      a => sym_counter_op_net_x0,
      b(0) => constant7_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  relational5: entity work.relational_9108cf519a
    port map (
      a => sym_counter_op_net_x0,
      b => constant8_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net
    );

  relational6: entity work.relational_9108cf519a
    port map (
      a => sym_counter_op_net_x0,
      b => constant9_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational6_op_net
    );

  relational7: entity work.relational_5b4e5df320
    port map (
      a => sym_counter_op_net_x0,
      b => constant10_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational7_op_net
    );

  x2lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 10,
      y_width => 2
    )
    port map (
      x => sym_counter_op_net_x0,
      y => x2lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/OFDM Symbol Ctrl/Sym Counter"

entity sym_counter_entity_fb3e36dd76 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    start_sym: in std_logic; 
    tx_reset: in std_logic; 
    start_sym_x0: out std_logic; 
    sym_ind: out std_logic_vector(9 downto 0)
  );
end sym_counter_entity_fb3e36dd76;

architecture structural of sym_counter_entity_fb3e36dd76 is
  signal ce_1_sg_x16: std_logic;
  signal clk_1_sg_x16: std_logic;
  signal delay_q_net_x0: std_logic;
  signal logical2_y_net: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net_x8: std_logic;
  signal register2_q_net_x0: std_logic;
  signal sym_counter_op_net_x1: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x16 <= ce_1;
  clk_1_sg_x16 <= clk_1;
  logical2_y_net_x1 <= start_sym;
  logical_y_net_x8 <= tx_reset;
  start_sym_x0 <= delay_q_net_x0;
  sym_ind <= sym_counter_op_net_x1;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      d(0) => logical2_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x0
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical2_y_net_x1,
      d1(0) => register2_q_net_x0,
      y(0) => logical2_y_net
    );

  s_r_latch1_b6e3de9a37: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x16,
      clk_1 => clk_1_sg_x16,
      r => logical_y_net_x8,
      s => logical2_y_net_x1,
      q => register2_q_net_x0
    );

  sym_counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      clr => '0',
      en(0) => logical2_y_net,
      rst(0) => logical_y_net_x8,
      op => sym_counter_op_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/OFDM Symbol Ctrl/Sym Samp Counter"

entity sym_samp_counter_entity_a7b82cdcb9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    sym_cfg: in std_logic_vector(17 downto 0); 
    sym_started: in std_logic; 
    tx_iq_samp_ce: in std_logic; 
    tx_reset: in std_logic; 
    start_next: out std_logic
  );
end sym_samp_counter_entity_a7b82cdcb9;

architecture structural of sym_samp_counter_entity_a7b82cdcb9 is
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal ce_1_sg_x20: std_logic;
  signal clk_1_sg_x20: std_logic;
  signal concat_y_net_x3: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical2_y_net: std_logic;
  signal logical4_y_net_x3: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x9: std_logic;
  signal mcode_cyclic_prefix_net: std_logic_vector(4 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register8_q_net_x3: std_logic_vector(7 downto 0);
  signal relational2_op_net_x0: std_logic;
  signal samp_counter_op_net: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x20 <= ce_1;
  clk_1_sg_x20 <= clk_1;
  register8_q_net_x3 <= regtx_num_sc;
  concat_y_net_x3 <= sym_cfg;
  logical4_y_net_x3 <= sym_started;
  convert2_dout_net_x0 <= tx_iq_samp_ce;
  logical_y_net_x9 <= tx_reset;
  start_next <= logical1_y_net_x3;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 5,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 9,
      core_name0 => "addsb_11_0_60fd3b5996582b7a",
      en_arith => xlUnsigned,
      en_bin_pt => 0,
      en_width => 1,
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 9,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => register8_q_net_x3,
      b => mcode_cyclic_prefix_net,
      ce => ce_1_sg_x20,
      clk => clk_1_sg_x20,
      clr => '0',
      en(0) => logical_y_net_x9,
      s => addsub_s_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x20,
      clk => clk_1_sg_x20,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => convert2_dout_net_x0,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x9,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x9,
      d1(0) => inverter_op_net,
      y(0) => logical2_y_net
    );

  mcode: entity work.mcode_block_00412594a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      sym_cfg => concat_y_net_x3,
      cyclic_prefix => mcode_cyclic_prefix_net
    );

  posedge1_e2905cab04: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x20,
      clk_1 => clk_1_sg_x20,
      d => logical4_y_net_x3,
      q => logical1_y_net_x2
    );

  posedge2_fd3e7298ed: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x20,
      clk_1 => clk_1_sg_x20,
      d => relational2_op_net_x0,
      q => logical1_y_net_x3
    );

  relational2: entity work.relational_6158158994
    port map (
      a => samp_counter_op_net,
      b => addsub_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net_x0
    );

  s_r_latch2_810e88f8a9: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x20,
      clk_1 => clk_1_sg_x20,
      r => logical1_y_net_x1,
      s => logical1_y_net_x2,
      q => register2_q_net_x0
    );

  samp_counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x20,
      clk => clk_1_sg_x20,
      clr => '0',
      en(0) => logical_y_net,
      rst(0) => logical2_y_net,
      op => samp_counter_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/OFDM Symbol Ctrl"

entity ofdm_symbol_ctrl_entity_c16241a486 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    convert2: in std_logic; 
    data_done: in std_logic; 
    logical3_x0: in std_logic; 
    output_fifo_occ: in std_logic_vector(7 downto 0); 
    register8: in std_logic_vector(7 downto 0); 
    slice: in std_logic; 
    slice1: in std_logic; 
    start_tx: in std_logic; 
    sym_done: in std_logic; 
    tx_reset: in std_logic; 
    start_sym: out std_logic; 
    sym_cfg: out std_logic_vector(17 downto 0)
  );
end ofdm_symbol_ctrl_entity_c16241a486;

architecture structural of ofdm_symbol_ctrl_entity_c16241a486 is
  signal ce_1_sg_x21: std_logic;
  signal clk_1_sg_x21: std_logic;
  signal concat_y_net_x4: std_logic_vector(17 downto 0);
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal convert2_dout_net_x1: std_logic;
  signal delay9_q_net_x1: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fifo_dcount_net_x0: std_logic_vector(7 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical3_y_net: std_logic;
  signal logical3_y_net_x2: std_logic;
  signal logical4_y_net_x4: std_logic;
  signal logical5_y_net: std_logic;
  signal logical_y_net_x10: std_logic;
  signal mux3_y_net_x3: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x2: std_logic;
  signal register3_q_net_x1: std_logic;
  signal register8_q_net_x4: std_logic_vector(7 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net_x0: std_logic;
  signal slice1_y_net_x1: std_logic;
  signal slice_y_net_x1: std_logic;
  signal sym_counter_op_net_x1: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x21 <= ce_1;
  clk_1_sg_x21 <= clk_1;
  convert2_dout_net_x1 <= convert2;
  delay9_q_net_x1 <= data_done;
  logical3_y_net_x2 <= logical3_x0;
  fifo_dcount_net_x0 <= output_fifo_occ;
  register8_q_net_x4 <= register8;
  slice_y_net_x1 <= slice;
  slice1_y_net_x1 <= slice1;
  register3_q_net_x1 <= start_tx;
  mux3_y_net_x3 <= sym_done;
  logical_y_net_x10 <= tx_reset;
  start_sym <= logical4_y_net_x4;
  sym_cfg <= concat_y_net_x4;

  constant1: entity work.constant_b8fb990c43
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x21,
      clk => clk_1_sg_x21,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x21,
      clk => clk_1_sg_x21,
      clr => '0',
      ip(0) => register2_q_net_x2,
      op(0) => inverter2_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x2,
      d1(0) => logical1_y_net_x4,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_a6d07705dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => logical3_y_net,
      d2(0) => logical5_y_net,
      d3(0) => logical1_y_net,
      y(0) => logical2_y_net_x1
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net,
      d1(0) => mux3_y_net_x3,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => inverter1_op_net,
      d2(0) => register2_q_net_x1,
      y(0) => logical4_y_net_x4
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x2,
      d1(0) => inverter2_op_net,
      y(0) => logical5_y_net
    );

  posedge1_78541e5bea: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      d => register3_q_net_x1,
      q => logical1_y_net_x1
    );

  posedge2_9f3bdafa2c: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      d => relational2_op_net_x0,
      q => logical1_y_net_x2
    );

  posedge3_2b1b2320ea: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      d => delay9_q_net_x1,
      q => logical1_y_net_x3
    );

  relational1: entity work.relational_ecce2f20df
    port map (
      a => sym_counter_op_net_x1,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_2d417722ee
    port map (
      a => fifo_dcount_net_x0,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net_x0
    );

  s_r_latch1_04de4f2c71: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      r => logical_y_net_x10,
      s => logical1_y_net_x3,
      q => register2_q_net_x0
    );

  s_r_latch2_7f5a15fb9e: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      r => logical_y_net_x10,
      s => logical1_y_net_x1,
      q => register2_q_net_x1
    );

  s_r_latch3_08b9ae30e7: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      r => logical_y_net_x10,
      s => logical1_y_net_x2,
      q => register2_q_net_x2
    );

  sym_config_encode_43a940459d: entity work.sym_config_encode_entity_43a940459d
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      ofdm_sym_ind => sym_counter_op_net_x1,
      tx_phy_mode_11ag => slice_y_net_x1,
      tx_phy_mode_11n => slice1_y_net_x1,
      tx_phy_mode_11n_ac => logical3_y_net_x2,
      sym_cfg => concat_y_net_x4
    );

  sym_counter_fb3e36dd76: entity work.sym_counter_entity_fb3e36dd76
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      start_sym => logical2_y_net_x1,
      tx_reset => logical_y_net_x10,
      start_sym_x0 => delay_q_net_x0,
      sym_ind => sym_counter_op_net_x1
    );

  sym_samp_counter_a7b82cdcb9: entity work.sym_samp_counter_entity_a7b82cdcb9
    port map (
      ce_1 => ce_1_sg_x21,
      clk_1 => clk_1_sg_x21,
      regtx_num_sc => register8_q_net_x4,
      sym_cfg => concat_y_net_x4,
      sym_started => logical4_y_net_x4,
      tx_iq_samp_ce => convert2_dout_net_x1,
      tx_reset => logical_y_net_x10,
      start_next => logical1_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Convolutional Encoder"

entity convolutional_encoder_entity_c777b8e511 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    tx_bit: in std_logic; 
    tx_bit_tlast: in std_logic; 
    tx_bit_tvalid: in std_logic; 
    tx_reset: in std_logic; 
    enc_bit_a: out std_logic; 
    enc_bit_b: out std_logic; 
    enc_bits_tlast: out std_logic; 
    enc_bits_tvalid: out std_logic; 
    sym_cfg_x0: out std_logic_vector(17 downto 0)
  );
end convolutional_encoder_entity_c777b8e511;

architecture structural of convolutional_encoder_entity_c777b8e511 is
  signal a_xor_y_net_x0: std_logic;
  signal b_xor_y_net_x0: std_logic;
  signal ce_1_sg_x22: std_logic;
  signal clk_1_sg_x22: std_logic;
  signal convert2_dout_net: std_logic;
  signal convert_dout_net: std_logic;
  signal delay1_q_net_x0: std_logic_vector(17 downto 0);
  signal delay2_q_net_x1: std_logic;
  signal delay2_q_net_x2: std_logic;
  signal delay3_q_net_x0: std_logic;
  signal delay8_q_net_x0: std_logic_vector(17 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x11: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x22 <= ce_1;
  clk_1_sg_x22 <= clk_1;
  delay8_q_net_x0 <= sym_cfg;
  logical_y_net_x0 <= tx_bit;
  logical1_y_net_x0 <= tx_bit_tlast;
  delay2_q_net_x1 <= tx_bit_tvalid;
  logical_y_net_x11 <= tx_reset;
  enc_bit_a <= a_xor_y_net_x0;
  enc_bit_b <= b_xor_y_net_x0;
  enc_bits_tlast <= delay2_q_net_x2;
  enc_bits_tvalid <= delay3_q_net_x0;
  sym_cfg_x0 <= delay1_q_net_x0;

  a_xor: entity work.logical_899cf9b568
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      d0(0) => logical_y_net_x0,
      d1(0) => register1_q_net,
      d2(0) => register2_q_net,
      d3(0) => register4_q_net,
      d4(0) => register5_q_net,
      en(0) => convert2_dout_net,
      y(0) => a_xor_y_net_x0
    );

  b_xor: entity work.logical_899cf9b568
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      d0(0) => logical_y_net_x0,
      d1(0) => register_q_net,
      d2(0) => register1_q_net,
      d3(0) => register2_q_net,
      d4(0) => register5_q_net,
      en(0) => convert2_dout_net,
      y(0) => b_xor_y_net_x0
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      din(0) => logical_y_net_x11,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      din(0) => delay2_q_net_x1,
      en => "1",
      dout(0) => convert2_dout_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d => delay8_q_net_x0,
      en => '1',
      rst => '1',
      q => delay1_q_net_x0
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => logical1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x2
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => convert2_dout_net,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => register_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => register1_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => register2_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => register3_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => register4_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      d(0) => logical_y_net_x0,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Index Gen/Bit Index Gen"

entity bit_index_gen_entity_9506081c38 is
  port (
    bit_rd_en: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    tx_reset: in std_logic; 
    bit_sel: out std_logic_vector(2 downto 0); 
    byte_ind: out std_logic_vector(11 downto 0); 
    byte_ind_valid: out std_logic
  );
end bit_index_gen_entity_9506081c38;

architecture structural of bit_index_gen_entity_9506081c38 is
  signal bit_counter_op_net: std_logic_vector(14 downto 0);
  signal bit_in_byte_y_net_x0: std_logic_vector(2 downto 0);
  signal bytes_y_net_x0: std_logic_vector(11 downto 0);
  signal ce_1_sg_x23: std_logic;
  signal clk_1_sg_x23: std_logic;
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal logical4_y_net_x0: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net_x12: std_logic;
  signal relational1_op_net: std_logic;

begin
  logical4_y_net_x0 <= bit_rd_en;
  ce_1_sg_x23 <= ce_1;
  clk_1_sg_x23 <= clk_1;
  logical_y_net_x12 <= tx_reset;
  bit_sel <= bit_in_byte_y_net_x0;
  byte_ind <= bytes_y_net_x0;
  byte_ind_valid <= logical5_y_net_x0;

  bit_counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_d5912692bc2e79ac",
      op_arith => xlUnsigned,
      op_width => 15
    )
    port map (
      ce => ce_1_sg_x23,
      clk => clk_1_sg_x23,
      clr => '0',
      en(0) => logical4_y_net_x0,
      rst(0) => logical_y_net_x12,
      op => bit_counter_op_net
    );

  bit_in_byte: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 15,
      y_width => 3
    )
    port map (
      x => bit_counter_op_net,
      y => bit_in_byte_y_net_x0
    );

  bytes: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 14,
      x_width => 15,
      y_width => 12
    )
    port map (
      x => bit_counter_op_net,
      y => bytes_y_net_x0
    );

  constant3: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net,
      d1(0) => logical4_y_net_x0,
      y(0) => logical5_y_net_x0
    );

  relational1: entity work.relational_706b9eb7ce
    port map (
      a => bit_in_byte_y_net_x0,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Index Gen/Bits Per Sym"

entity bits_per_sym_entity_70418c6109 is
  port (
    base_rate: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    full_rate: in std_logic; 
    ofdm_tx_data_n_dbps: in std_logic_vector(9 downto 0); 
    start: in std_logic; 
    tx_reset: in std_logic; 
    rd_en: out std_logic
  );
end bits_per_sym_entity_70418c6109;

architecture structural of bits_per_sym_entity_70418c6109 is
  signal ce_1_sg_x25: std_logic;
  signal clk_1_sg_x25: std_logic;
  signal constant2_op_net: std_logic_vector(4 downto 0);
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical4_y_net_x1: std_logic;
  signal logical4_y_net_x5: std_logic;
  signal logical_y_net_x13: std_logic;
  signal mcode_load_base_rate_net_x0: std_logic;
  signal mcode_load_full_rate_net_x0: std_logic;
  signal mux_y_net: std_logic_vector(9 downto 0);
  signal register1_q_net_x0: std_logic_vector(9 downto 0);
  signal register2_q_net: std_logic_vector(9 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register3_q_net: std_logic;
  signal relational3_op_net: std_logic;

begin
  mcode_load_base_rate_net_x0 <= base_rate;
  ce_1_sg_x25 <= ce_1;
  clk_1_sg_x25 <= clk_1;
  mcode_load_full_rate_net_x0 <= full_rate;
  register1_q_net_x0 <= ofdm_tx_data_n_dbps;
  logical4_y_net_x5 <= start;
  logical_y_net_x13 <= tx_reset;
  rd_en <= logical4_y_net_x1;

  constant2: entity work.constant_bc74ae1a6c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      clr => '0',
      en(0) => register2_q_net_x0,
      rst(0) => inverter1_op_net,
      op => counter_op_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      clr => '0',
      ip(0) => relational3_op_net,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x13,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net_x0
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => mcode_load_full_rate_net_x0,
      d1(0) => mcode_load_base_rate_net_x0,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical4_y_net_x5,
      d1(0) => logical2_y_net,
      y(0) => logical3_y_net_x0
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => register2_q_net_x0,
      y(0) => logical4_y_net_x1
    );

  mux: entity work.mux_02d5ef99fc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register2_q_net,
      d1 => constant2_op_net,
      sel(0) => register3_q_net,
      y => mux_y_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 10,
      init_value => b"0000011000"
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d => register1_q_net_x0,
      en(0) => logical3_y_net_x0,
      rst(0) => logical_y_net_x13,
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => mcode_load_base_rate_net_x0,
      en(0) => logical3_y_net_x0,
      rst(0) => logical_y_net_x13,
      q(0) => register3_q_net
    );

  relational3: entity work.relational_1813613113
    port map (
      a => counter_op_net,
      b => mux_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_696cea2643: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      r => logical1_y_net_x0,
      s => logical3_y_net_x0,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Index Gen"

entity index_gen_entity_b965cbdf90 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    logical: in std_logic; 
    register1: in std_logic_vector(9 downto 0); 
    start_sym: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    bit_sel: out std_logic_vector(2 downto 0); 
    bit_sel_valid: out std_logic; 
    byte_ind: out std_logic_vector(11 downto 0); 
    byte_ind_valid: out std_logic
  );
end index_gen_entity_b965cbdf90;

architecture structural of index_gen_entity_b965cbdf90 is
  signal bit_in_byte_y_net_x1: std_logic_vector(2 downto 0);
  signal bytes_y_net_x1: std_logic_vector(11 downto 0);
  signal ce_1_sg_x26: std_logic;
  signal clk_1_sg_x26: std_logic;
  signal concat_y_net_x5: std_logic_vector(17 downto 0);
  signal logical4_y_net_x2: std_logic;
  signal logical4_y_net_x6: std_logic;
  signal logical5_y_net_x1: std_logic;
  signal logical_y_net_x14: std_logic;
  signal mcode_load_base_rate_net_x0: std_logic;
  signal mcode_load_full_rate_net_x0: std_logic;
  signal register1_q_net_x1: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x26 <= ce_1;
  clk_1_sg_x26 <= clk_1;
  logical_y_net_x14 <= logical;
  register1_q_net_x1 <= register1;
  logical4_y_net_x6 <= start_sym;
  concat_y_net_x5 <= sym_cfg;
  bit_sel <= bit_in_byte_y_net_x1;
  bit_sel_valid <= logical4_y_net_x2;
  byte_ind <= bytes_y_net_x1;
  byte_ind_valid <= logical5_y_net_x1;

  bit_index_gen_9506081c38: entity work.bit_index_gen_entity_9506081c38
    port map (
      bit_rd_en => logical4_y_net_x2,
      ce_1 => ce_1_sg_x26,
      clk_1 => clk_1_sg_x26,
      tx_reset => logical_y_net_x14,
      bit_sel => bit_in_byte_y_net_x1,
      byte_ind => bytes_y_net_x1,
      byte_ind_valid => logical5_y_net_x1
    );

  bits_per_sym_70418c6109: entity work.bits_per_sym_entity_70418c6109
    port map (
      base_rate => mcode_load_base_rate_net_x0,
      ce_1 => ce_1_sg_x26,
      clk_1 => clk_1_sg_x26,
      full_rate => mcode_load_full_rate_net_x0,
      ofdm_tx_data_n_dbps => register1_q_net_x1,
      start => logical4_y_net_x6,
      tx_reset => logical_y_net_x14,
      rd_en => logical4_y_net_x2
    );

  mcode: entity work.mcode_block_00412594a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      sym_cfg => concat_y_net_x5,
      load_base_rate(0) => mcode_load_base_rate_net_x0,
      load_full_rate(0) => mcode_load_full_rate_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/16QAM Mod"

entity x16qam_mod_entity_19a899dd5b is
  port (
    b_3_0: in std_logic_vector(3 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end x16qam_mod_entity_19a899dd5b;

architecture structural of x16qam_mod_entity_19a899dd5b is
  signal b_1_0_y_net: std_logic_vector(1 downto 0);
  signal b_3_2_y_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal x4lsb_y_net_x0: std_logic_vector(3 downto 0);

begin
  x4lsb_y_net_x0 <= b_3_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  b_1_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => x4lsb_y_net_x0,
      y => b_1_0_y_net
    );

  b_3_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => x4lsb_y_net_x0,
      y => b_3_2_y_net
    );

  constant1: entity work.constant_fd8727242d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_c09b53cba3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_41d1fb8f4c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_aec943c743
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  mux: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      sel => b_1_0_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      sel => b_3_2_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/64QAM Mod"

entity x64qam_mod_entity_51e5e09af7 is
  port (
    b_5_0: in std_logic_vector(5 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end x64qam_mod_entity_51e5e09af7;

architecture structural of x64qam_mod_entity_51e5e09af7 is
  signal b_2_0_y_net: std_logic_vector(2 downto 0);
  signal b_5_3_y_net: std_logic_vector(2 downto 0);
  signal constant10_op_net: std_logic_vector(11 downto 0);
  signal constant11_op_net: std_logic_vector(11 downto 0);
  signal constant12_op_net: std_logic_vector(11 downto 0);
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal constant9_op_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal x6lsb_y_net_x0: std_logic_vector(5 downto 0);

begin
  x6lsb_y_net_x0 <= b_5_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  b_2_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 6,
      y_width => 3
    )
    port map (
      x => x6lsb_y_net_x0,
      y => b_2_0_y_net
    );

  b_5_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 5,
      x_width => 6,
      y_width => 3
    )
    port map (
      x => x6lsb_y_net_x0,
      y => b_5_3_y_net
    );

  constant1: entity work.constant_9127ce6619
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant10: entity work.constant_50239c0b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant10_op_net
    );

  constant11: entity work.constant_1971ed2879
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant11_op_net
    );

  constant12: entity work.constant_93635891b9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant12_op_net
    );

  constant2: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_9fcec64691
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_8da791e271
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant9: entity work.constant_c3ad5f20a9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant9_op_net
    );

  mux: entity work.mux_f3bb14635d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      d4 => constant10_op_net,
      d5 => constant9_op_net,
      d6 => constant11_op_net,
      d7 => constant12_op_net,
      sel => b_2_0_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_f3bb14635d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      d4 => constant10_op_net,
      d5 => constant9_op_net,
      d6 => constant11_op_net,
      d7 => constant12_op_net,
      sel => b_5_3_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/BPSK Mod"

entity bpsk_mod_entity_12640088e5 is
  port (
    b_0: in std_logic; 
    rot: in std_logic; 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end bpsk_mod_entity_12640088e5;

architecture structural of bpsk_mod_entity_12640088e5 is
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal mcode_rotate_bpsk_net_x0: std_logic;
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux2_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal x1lsb_y_net_x0: std_logic;

begin
  x1lsb_y_net_x0 <= b_0;
  mcode_rotate_bpsk_net_x0 <= rot;
  i <= mux1_y_net_x0;
  q <= mux2_y_net_x0;

  constant2: entity work.constant_7e4d1a10e6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_afc893bf70
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  mux: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => x1lsb_y_net_x0,
      y => mux_y_net
    );

  mux1: entity work.mux_4de2214a42
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux_y_net,
      d1 => constant4_op_net,
      sel(0) => mcode_rotate_bpsk_net_x0,
      y => mux1_y_net_x0
    );

  mux2: entity work.mux_4de2214a42
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant4_op_net,
      d1 => mux_y_net,
      sel(0) => mcode_rotate_bpsk_net_x0,
      y => mux2_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots/Data SC Map"

entity data_sc_map_entity_45d00f2f68 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    full_rate: in std_logic; 
    sc_ind: in std_logic_vector(5 downto 0); 
    tx_phy_mode_11n: in std_logic; 
    data_sym_ind: out std_logic_vector(5 downto 0); 
    data_sym_valid: out std_logic
  );
end data_sc_map_entity_45d00f2f68;

architecture structural of data_sc_map_entity_45d00f2f68 is
  signal ce_1_sg_x27: std_logic;
  signal clk_1_sg_x27: std_logic;
  signal constant2_op_net: std_logic_vector(6 downto 0);
  signal logical_y_net: std_logic;
  signal mcode_load_full_rate_net_x0: std_logic;
  signal mux1_y_net: std_logic_vector(6 downto 0);
  signal relational1_op_net_x0: std_logic;
  signal slice1_y_net_x2: std_logic;
  signal slice_y_net_x0: std_logic_vector(5 downto 0);
  signal subcarrier_index_op_net_x0: std_logic_vector(5 downto 0);
  signal x11a_subcarrier_map_data_net: std_logic_vector(6 downto 0);
  signal x11n_ht20_subcarrier_map_data_net: std_logic_vector(6 downto 0);

begin
  ce_1_sg_x27 <= ce_1;
  clk_1_sg_x27 <= clk_1;
  mcode_load_full_rate_net_x0 <= full_rate;
  subcarrier_index_op_net_x0 <= sc_ind;
  slice1_y_net_x2 <= tx_phy_mode_11n;
  data_sym_ind <= slice_y_net_x0;
  data_sym_valid <= relational1_op_net_x0;

  constant2: entity work.constant_7b07120b87
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x2,
      d1(0) => mcode_load_full_rate_net_x0,
      y(0) => logical_y_net
    );

  mux1: entity work.mux_3797c120ed
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => x11a_subcarrier_map_data_net,
      d1 => x11n_ht20_subcarrier_map_data_net,
      sel(0) => logical_y_net,
      y => mux1_y_net
    );

  relational1: entity work.relational_23065a6aa3
    port map (
      a => mux1_y_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 7,
      y_width => 6
    )
    port map (
      x => mux1_y_net,
      y => slice_y_net_x0
    );

  x11a_subcarrier_map: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 6,
      c_address_width => 6,
      c_width => 7,
      core_name0 => "dmg_72_58f1077b49388e77",
      latency => 0
    )
    port map (
      addr => subcarrier_index_op_net_x0,
      ce => ce_1_sg_x27,
      clk => clk_1_sg_x27,
      en => "1",
      data => x11a_subcarrier_map_data_net
    );

  x11n_ht20_subcarrier_map: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 6,
      c_address_width => 6,
      c_width => 7,
      core_name0 => "dmg_72_d59da422e431313e",
      latency => 0
    )
    port map (
      addr => subcarrier_index_op_net_x0,
      ce => ce_1_sg_x27,
      clk => clk_1_sg_x27,
      en => "1",
      data => x11n_ht20_subcarrier_map_data_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots/Pilot Gen/Pilot Selection"

entity pilot_selection_entity_35ea130450 is
  port (
    sc_ind: in std_logic_vector(5 downto 0); 
    shift: in std_logic_vector(1 downto 0); 
    negate: out std_logic; 
    pilot: out std_logic
  );
end pilot_selection_entity_35ea130450;

architecture structural of pilot_selection_entity_35ea130450 is
  signal constant1_op_net: std_logic_vector(5 downto 0);
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal constant3_op_net: std_logic_vector(5 downto 0);
  signal constant4_op_net: std_logic_vector(5 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal mcode_pilot_shift_net_x0: std_logic_vector(1 downto 0);
  signal mux_y_net_x0: std_logic;
  signal relational4_op_net: std_logic;
  signal relational5_op_net: std_logic;
  signal relational6_op_net: std_logic;
  signal relational7_op_net: std_logic;
  signal subcarrier_index_op_net_x1: std_logic_vector(5 downto 0);

begin
  subcarrier_index_op_net_x1 <= sc_ind;
  mcode_pilot_shift_net_x0 <= shift;
  negate <= mux_y_net_x0;
  pilot <= logical1_y_net_x0;

  constant1: entity work.constant_1f05b15a2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_330e503d71
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_173d83e4a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_8207020ee3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  logical1: entity work.logical_a6d07705dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational4_op_net,
      d1(0) => relational5_op_net,
      d2(0) => relational6_op_net,
      d3(0) => relational7_op_net,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_cdffdf53c9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational5_op_net,
      d1(0) => relational4_op_net,
      d2(0) => relational7_op_net,
      d3(0) => relational6_op_net,
      sel => mcode_pilot_shift_net_x0,
      y(0) => mux_y_net_x0
    );

  relational4: entity work.relational_931d61fb72
    port map (
      a => constant2_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  relational5: entity work.relational_931d61fb72
    port map (
      a => constant1_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net
    );

  relational6: entity work.relational_931d61fb72
    port map (
      a => constant4_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational6_op_net
    );

  relational7: entity work.relational_931d61fb72
    port map (
      a => constant3_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational7_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots/Pilot Gen/Scrambling LFSR"

entity scrambling_lfsr_entity_63498a346e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    q: out std_logic
  );
end scrambling_lfsr_entity_63498a346e;

architecture structural of scrambling_lfsr_entity_63498a346e is
  signal assert1_dout_net: std_logic;
  signal assert_dout_net: std_logic;
  signal ce_1_sg_x29: std_logic;
  signal clk_1_sg_x29: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x15: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register6_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x29 <= ce_1;
  clk_1_sg_x29 <= clk_1;
  logical1_y_net_x1 <= en;
  logical_y_net_x15 <= rst;
  q <= logical_y_net_x0;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register3_q_net,
      dout(0) => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register6_q_net,
      dout(0) => assert_dout_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din(0) => logical_y_net_x15,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din(0) => logical1_y_net_x1,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => assert_dout_net,
      d1(0) => assert1_dout_net,
      y(0) => logical_y_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register1_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register2_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register3_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register4_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => register5_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register6_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => logical_y_net_x0,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots/Pilot Gen"

entity pilot_gen_entity_da39436044 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    pilot_shift: in std_logic_vector(1 downto 0); 
    reset: in std_logic; 
    sc_ind: in std_logic_vector(5 downto 0); 
    pilot_i: out std_logic_vector(11 downto 0); 
    pilot_valid: out std_logic
  );
end pilot_gen_entity_da39436044;

architecture structural of pilot_gen_entity_da39436044 is
  signal ce_1_sg_x30: std_logic;
  signal clk_1_sg_x30: std_logic;
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant5_op_net: std_logic_vector(11 downto 0);
  signal delay_q_net: std_logic_vector(5 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x16: std_logic;
  signal mcode_pilot_shift_net_x1: std_logic_vector(1 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal subcarrier_index_op_net_x2: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x30 <= ce_1;
  clk_1_sg_x30 <= clk_1;
  mcode_pilot_shift_net_x1 <= pilot_shift;
  logical_y_net_x16 <= reset;
  subcarrier_index_op_net_x2 <= sc_ind;
  pilot_i <= mux1_y_net_x0;
  pilot_valid <= logical1_y_net_x2;

  constant1: entity work.constant_7e4d1a10e6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant5: entity work.constant_afc893bf70
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 6
    )
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      d => subcarrier_index_op_net_x2,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => mux_y_net_x0,
      d1(0) => logical_y_net_x0,
      y(0) => logical_y_net
    );

  mux1: entity work.mux_4de2214a42
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant5_op_net,
      d1 => constant1_op_net,
      sel(0) => logical_y_net,
      y => mux1_y_net_x0
    );

  pilot_selection_35ea130450: entity work.pilot_selection_entity_35ea130450
    port map (
      sc_ind => subcarrier_index_op_net_x2,
      shift => mcode_pilot_shift_net_x1,
      negate => mux_y_net_x0,
      pilot => logical1_y_net_x2
    );

  posedge_cc752e9a4c: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      d => relational1_op_net_x0,
      q => logical1_y_net_x1
    );

  relational1: entity work.relational_47932db5b1
    port map (
      a => subcarrier_index_op_net_x2,
      b => delay_q_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  scrambling_lfsr_63498a346e: entity work.scrambling_lfsr_entity_63498a346e
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      en => logical1_y_net_x1,
      rst => logical_y_net_x16,
      q => logical_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots/Subcarrier Index Count"

entity subcarrier_index_count_entity_37e2404044 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    reset: in std_logic; 
    last: out std_logic; 
    sc_ind: out std_logic_vector(5 downto 0)
  );
end subcarrier_index_count_entity_37e2404044;

architecture structural of subcarrier_index_count_entity_37e2404044 is
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal ce_1_sg_x34: std_logic;
  signal clk_1_sg_x34: std_logic;
  signal constant1_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net: std_logic;
  signal logical_y_net_x17: std_logic;
  signal register8_q_net_x5: std_logic_vector(7 downto 0);
  signal relational3_op_net: std_logic;
  signal subcarrier_index_op_net_x3: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x34 <= ce_1;
  clk_1_sg_x34 <= clk_1;
  logical1_y_net_x1 <= en;
  register8_q_net_x5 <= regtx_num_sc;
  logical_y_net_x17 <= reset;
  last <= logical1_y_net_x2;
  sc_ind <= subcarrier_index_op_net_x3;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 1,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 9,
      core_name0 => "addsb_11_0_a52ead9b8a3c1e76",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 9,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => register8_q_net_x5,
      b(0) => constant1_op_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x17,
      d1(0) => logical1_y_net_x2,
      y(0) => logical2_y_net
    );

  relational3: entity work.relational_1834ac00b4
    port map (
      a => addsub_s_net,
      b => subcarrier_index_op_net_x3,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  subcarrier_index: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_f068fb73312ae1e5",
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      en(0) => logical1_y_net_x1,
      rst(0) => logical2_y_net,
      op => subcarrier_index_op_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/Control & Pilots"

entity \control___pilots_entity_44c57f2255\ is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    full_rate: in std_logic; 
    iq_fifo_tready: in std_logic; 
    pilot_shift: in std_logic_vector(1 downto 0); 
    register8: in std_logic_vector(7 downto 0); 
    slice1: in std_logic; 
    sym_bits_rdy: in std_logic; 
    tx_reset: in std_logic; 
    data_sym_ind: out std_logic_vector(5 downto 0); 
    iq_sel: out std_logic_vector(1 downto 0); 
    iq_tlast: out std_logic; 
    iq_tvalid: out std_logic; 
    pilot_i: out std_logic_vector(11 downto 0)
  );
end \control___pilots_entity_44c57f2255\;

architecture structural of \control___pilots_entity_44c57f2255\ is
  signal axi_fifo_s_axis_tready_net_x3: std_logic;
  signal ce_1_sg_x35: std_logic;
  signal clk_1_sg_x35: std_logic;
  signal concat1_y_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x1: std_logic;
  signal delay5_q_net_x1: std_logic;
  signal delay5_q_net_x2: std_logic_vector(1 downto 0);
  signal delay6_q_net_x0: std_logic_vector(11 downto 0);
  signal delay_q_net_x4: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x18: std_logic;
  signal mcode_load_full_rate_net_x1: std_logic;
  signal mcode_pilot_shift_net_x2: std_logic_vector(1 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register8_q_net_x6: std_logic_vector(7 downto 0);
  signal relational1_op_net_x0: std_logic;
  signal slice1_y_net_x3: std_logic;
  signal slice_y_net_x1: std_logic_vector(5 downto 0);
  signal subcarrier_index_op_net_x3: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x35 <= ce_1;
  clk_1_sg_x35 <= clk_1;
  mcode_load_full_rate_net_x1 <= full_rate;
  axi_fifo_s_axis_tready_net_x3 <= iq_fifo_tready;
  mcode_pilot_shift_net_x2 <= pilot_shift;
  register8_q_net_x6 <= register8;
  slice1_y_net_x3 <= slice1;
  delay5_q_net_x1 <= sym_bits_rdy;
  logical_y_net_x18 <= tx_reset;
  data_sym_ind <= slice_y_net_x1;
  iq_sel <= delay5_q_net_x2;
  iq_tlast <= delay1_q_net_x1;
  iq_tvalid <= delay_q_net_x4;
  pilot_i <= delay6_q_net_x0;

  concat1: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => relational1_op_net_x0,
      in1(0) => logical1_y_net_x2,
      y => concat1_y_net
    );

  data_sc_map_45d00f2f68: entity work.data_sc_map_entity_45d00f2f68
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      full_rate => mcode_load_full_rate_net_x1,
      sc_ind => subcarrier_index_op_net_x3,
      tx_phy_mode_11n => slice1_y_net_x3,
      data_sym_ind => slice_y_net_x1,
      data_sym_valid => relational1_op_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x4
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d(0) => logical1_y_net_x5,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x1
    );

  delay5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 2
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => concat1_y_net,
      en => '1',
      rst => '1',
      q => delay5_q_net_x2
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => mux1_y_net_x0,
      en => '1',
      rst => '1',
      q => delay6_q_net_x0
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x18,
      d1(0) => logical1_y_net_x5,
      y(0) => logical_y_net_x0
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => axi_fifo_s_axis_tready_net_x3,
      y(0) => logical1_y_net_x1
    );

  pilot_gen_da39436044: entity work.pilot_gen_entity_da39436044
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      pilot_shift => mcode_pilot_shift_net_x2,
      reset => logical_y_net_x18,
      sc_ind => subcarrier_index_op_net_x3,
      pilot_i => mux1_y_net_x0,
      pilot_valid => logical1_y_net_x2
    );

  posedge1_7a697fced3: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      d => logical_y_net_x0,
      q => logical1_y_net_x4
    );

  posedge_fab6da5860: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      d => delay5_q_net_x1,
      q => logical1_y_net_x3
    );

  s_r_latch1_b90293cf40: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      r => logical1_y_net_x4,
      s => logical1_y_net_x3,
      q => register2_q_net_x0
    );

  subcarrier_index_count_37e2404044: entity work.subcarrier_index_count_entity_37e2404044
    port map (
      ce_1 => ce_1_sg_x35,
      clk_1 => clk_1_sg_x35,
      en => logical1_y_net_x1,
      regtx_num_sc => register8_q_net_x6,
      reset => logical_y_net_x18,
      last => logical1_y_net_x5,
      sc_ind => subcarrier_index_op_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate/QPSK Mod"

entity qpsk_mod_entity_7f9e653764 is
  port (
    b_1_0: in std_logic_vector(1 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end qpsk_mod_entity_7f9e653764;

architecture structural of qpsk_mod_entity_7f9e653764 is
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal lsb_1_y_net: std_logic;
  signal lsb_y_net: std_logic;
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal x2lsb_y_net_x0: std_logic_vector(1 downto 0);

begin
  x2lsb_y_net_x0 <= b_1_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  constant2: entity work.constant_cb767c7ef2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_d6a72b7a3b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => x2lsb_y_net_x0,
      y(0) => lsb_y_net
    );

  lsb_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => x2lsb_y_net_x0,
      y(0) => lsb_1_y_net
    );

  mux: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => lsb_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => lsb_1_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Modulate"

entity modulate_entity_324fd14050 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    iq_fifo_tready: in std_logic; 
    logical: in std_logic; 
    ofdm_tx_data_mod_sel: in std_logic_vector(1 downto 0); 
    register8: in std_logic_vector(7 downto 0); 
    sc_bits: in std_logic_vector(7 downto 0); 
    slice1: in std_logic; 
    sym_bits_rdy: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    data_sym_ind: out std_logic_vector(5 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    iq_tlast: out std_logic; 
    iq_tvalid: out std_logic; 
    q: out std_logic_vector(11 downto 0); 
    sym_cfg_x0: out std_logic_vector(17 downto 0)
  );
end modulate_entity_324fd14050;

architecture structural of modulate_entity_324fd14050 is
  signal axi_fifo_s_axis_tready_net_x4: std_logic;
  signal ce_1_sg_x36: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant5_op_net: std_logic_vector(11 downto 0);
  signal constant6_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x2: std_logic;
  signal delay5_q_net_x2: std_logic_vector(1 downto 0);
  signal delay5_q_net_x3: std_logic;
  signal delay6_q_net_x0: std_logic_vector(11 downto 0);
  signal delay6_q_net_x1: std_logic_vector(17 downto 0);
  signal delay_q_net_x6: std_logic;
  signal delay_q_net_x7: std_logic_vector(17 downto 0);
  signal logical2_y_net: std_logic_vector(1 downto 0);
  signal logical_y_net_x19: std_logic;
  signal mcode_load_full_rate_net_x1: std_logic;
  signal mcode_pilot_shift_net_x2: std_logic_vector(1 downto 0);
  signal mcode_rotate_bpsk_net_x0: std_logic;
  signal mux1_y_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux1_y_net_x1: std_logic_vector(11 downto 0);
  signal mux1_y_net_x2: std_logic_vector(11 downto 0);
  signal mux1_y_net_x3: std_logic_vector(11 downto 0);
  signal mux1_y_net_x5: std_logic_vector(7 downto 0);
  signal mux2_y_net: std_logic_vector(11 downto 0);
  signal mux2_y_net_x0: std_logic_vector(11 downto 0);
  signal mux3_y_net_x1: std_logic_vector(11 downto 0);
  signal mux4_y_net_x1: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x1: std_logic_vector(11 downto 0);
  signal mux_y_net_x2: std_logic_vector(11 downto 0);
  signal register2_q_net_x0: std_logic_vector(1 downto 0);
  signal register8_q_net_x7: std_logic_vector(7 downto 0);
  signal slice1_y_net_x4: std_logic;
  signal slice_y_net_x2: std_logic_vector(5 downto 0);
  signal x1lsb_y_net_x0: std_logic;
  signal x2lsb_y_net_x0: std_logic_vector(1 downto 0);
  signal x4lsb_y_net_x0: std_logic_vector(3 downto 0);
  signal x6lsb_y_net_x0: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x36 <= ce_1;
  clk_1_sg_x36 <= clk_1;
  axi_fifo_s_axis_tready_net_x4 <= iq_fifo_tready;
  logical_y_net_x19 <= logical;
  register2_q_net_x0 <= ofdm_tx_data_mod_sel;
  register8_q_net_x7 <= register8;
  mux1_y_net_x5 <= sc_bits;
  slice1_y_net_x4 <= slice1;
  delay5_q_net_x3 <= sym_bits_rdy;
  delay6_q_net_x1 <= sym_cfg;
  data_sym_ind <= slice_y_net_x2;
  i <= mux3_y_net_x1;
  iq_tlast <= delay1_q_net_x2;
  iq_tvalid <= delay_q_net_x6;
  q <= mux4_y_net_x1;
  sym_cfg_x0 <= delay_q_net_x7;

  bpsk_mod_12640088e5: entity work.bpsk_mod_entity_12640088e5
    port map (
      b_0 => x1lsb_y_net_x0,
      rot => mcode_rotate_bpsk_net_x0,
      i => mux1_y_net_x2,
      q => mux2_y_net_x0
    );

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => mcode_load_full_rate_net_x1,
      in1(0) => mcode_load_full_rate_net_x1,
      y => concat_y_net
    );

  constant5: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  control_pilots_44c57f2255: entity work.\control___pilots_entity_44c57f2255\
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      full_rate => mcode_load_full_rate_net_x1,
      iq_fifo_tready => axi_fifo_s_axis_tready_net_x4,
      pilot_shift => mcode_pilot_shift_net_x2,
      register8 => register8_q_net_x7,
      slice1 => slice1_y_net_x4,
      sym_bits_rdy => delay5_q_net_x3,
      tx_reset => logical_y_net_x19,
      data_sym_ind => slice_y_net_x2,
      iq_sel => delay5_q_net_x2,
      iq_tlast => delay1_q_net_x2,
      iq_tvalid => delay_q_net_x6,
      pilot_i => delay6_q_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d => delay6_q_net_x1,
      en => '1',
      rst => '1',
      q => delay_q_net_x7
    );

  logical2: entity work.logical_33c9a0c803
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat_y_net,
      d1 => register2_q_net_x0,
      y => logical2_y_net
    );

  mcode: entity work.mcode_block_00412594a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      sym_cfg => delay6_q_net_x1,
      load_full_rate(0) => mcode_load_full_rate_net_x1,
      pilot_shift => mcode_pilot_shift_net_x2,
      rotate_bpsk(0) => mcode_rotate_bpsk_net_x0
    );

  mux1: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux1_y_net_x2,
      d1 => mux_y_net_x2,
      d2 => mux_y_net_x0,
      d3 => mux_y_net_x1,
      sel => logical2_y_net,
      y => mux1_y_net
    );

  mux2: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux2_y_net_x0,
      d1 => mux1_y_net_x3,
      d2 => mux1_y_net_x0,
      d3 => mux1_y_net_x1,
      sel => logical2_y_net,
      y => mux2_y_net
    );

  mux3: entity work.mux_e5a9964709
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant6_op_net,
      d1 => delay6_q_net_x0,
      d2 => mux1_y_net,
      sel => delay5_q_net_x2,
      y => mux3_y_net_x1
    );

  mux4: entity work.mux_e5a9964709
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant5_op_net,
      d1 => constant5_op_net,
      d2 => mux2_y_net,
      sel => delay5_q_net_x2,
      y => mux4_y_net_x1
    );

  qpsk_mod_7f9e653764: entity work.qpsk_mod_entity_7f9e653764
    port map (
      b_1_0 => x2lsb_y_net_x0,
      i => mux_y_net_x2,
      q => mux1_y_net_x3
    );

  x16qam_mod_19a899dd5b: entity work.x16qam_mod_entity_19a899dd5b
    port map (
      b_3_0 => x4lsb_y_net_x0,
      i => mux_y_net_x0,
      q => mux1_y_net_x0
    );

  x1lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x5,
      y(0) => x1lsb_y_net_x0
    );

  x2lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => mux1_y_net_x5,
      y => x2lsb_y_net_x0
    );

  x4lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 8,
      y_width => 4
    )
    port map (
      x => mux1_y_net_x5,
      y => x4lsb_y_net_x0
    );

  x64qam_mod_51e5e09af7: entity work.x64qam_mod_entity_51e5e09af7
    port map (
      b_5_0 => x6lsb_y_net_x0,
      i => mux_y_net_x1,
      q => mux1_y_net_x1
    );

  x6lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => mux1_y_net_x5,
      y => x6lsb_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/BRAM IF 64b/BRAM Addr Map"

entity bram_addr_map_entity_8b602ce2fb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    tx_ind: in std_logic_vector(11 downto 0); 
    tx_phy_mode_11n_ac: in std_logic; 
    mem_addr: out std_logic_vector(11 downto 0)
  );
end bram_addr_map_entity_8b602ce2fb;

architecture structural of bram_addr_map_entity_8b602ce2fb is
  signal addsub1_s_net: std_logic_vector(11 downto 0);
  signal ce_1_sg_x37: std_logic;
  signal clk_1_sg_x37: std_logic;
  signal constant1_op_net: std_logic_vector(2 downto 0);
  signal constant2_op_net: std_logic_vector(3 downto 0);
  signal constant3_op_net: std_logic_vector(3 downto 0);
  signal constant4_op_net: std_logic_vector(2 downto 0);
  signal logical3_y_net_x3: std_logic;
  signal mux1_y_net: std_logic_vector(3 downto 0);
  signal mux2_y_net: std_logic_vector(3 downto 0);
  signal mux5_y_net_x0: std_logic_vector(11 downto 0);
  signal relational_op_net: std_logic;
  signal x12_lsb_y_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x37 <= ce_1;
  clk_1_sg_x37 <= clk_1;
  x12_lsb_y_net_x0 <= tx_ind;
  logical3_y_net_x3 <= tx_phy_mode_11n_ac;
  mem_addr <= mux5_y_net_x0;

  addsub1: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 12,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 4,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 13,
      core_name0 => "addsb_11_0_7cf14debcedb76ce",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 13,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 12
    )
    port map (
      a => x12_lsb_y_net_x0,
      b => mux2_y_net,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      clr => '0',
      en => "1",
      s => addsub1_s_net
    );

  constant1: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_c0ce4ae10c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_5c1626e05e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  mux1: entity work.mux_1e60cf48bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant1_op_net,
      d1 => constant3_op_net,
      sel(0) => logical3_y_net_x3,
      y => mux1_y_net
    );

  mux2: entity work.mux_102f86419c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant4_op_net,
      sel(0) => logical3_y_net_x3,
      y => mux2_y_net
    );

  mux5: entity work.mux_4de2214a42
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => addsub1_s_net,
      d1 => x12_lsb_y_net_x0,
      sel(0) => relational_op_net,
      y => mux5_y_net_x0
    );

  relational: entity work.relational_b218b04ee6
    port map (
      a => x12_lsb_y_net_x0,
      b => mux1_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/BRAM IF 64b/BRAM Interface"

entity bram_interface_entity_5cb2ccffdd is
  port (
    bram_din: in std_logic_vector(63 downto 0); 
    pkt_buf_index: in std_logic_vector(3 downto 0); 
    x64b_word_addr: in std_logic_vector(8 downto 0); 
    concat_x0: out std_logic_vector(31 downto 0); 
    constant1_x0: out std_logic; 
    constant2_x0: out std_logic; 
    constant7_x0: out std_logic_vector(63 downto 0); 
    constant8_x0: out std_logic_vector(7 downto 0); 
    x64b_data: out std_logic_vector(63 downto 0)
  );
end bram_interface_entity_5cb2ccffdd;

architecture structural of bram_interface_entity_5cb2ccffdd is
  signal addsub_s_net_x0: std_logic_vector(8 downto 0);
  signal bram_din_net_x0: std_logic_vector(63 downto 0);
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant1_op_net_x0: std_logic;
  signal constant2_op_net_x0: std_logic;
  signal constant3_op_net: std_logic_vector(2 downto 0);
  signal constant4_op_net: std_logic_vector(15 downto 0);
  signal constant7_op_net_x0: std_logic_vector(63 downto 0);
  signal constant8_op_net_x0: std_logic_vector(7 downto 0);
  signal mux_y_net_x0: std_logic_vector(3 downto 0);
  signal simulation_multiplexer_dout_net_x0: std_logic_vector(63 downto 0);

begin
  bram_din_net_x0 <= bram_din;
  mux_y_net_x0 <= pkt_buf_index;
  addsub_s_net_x0 <= x64b_word_addr;
  concat_x0 <= concat_y_net_x0;
  constant1_x0 <= constant1_op_net_x0;
  constant2_x0 <= constant2_op_net_x0;
  constant7_x0 <= constant7_op_net_x0;
  constant8_x0 <= constant8_op_net_x0;
  x64b_data <= simulation_multiplexer_dout_net_x0;

  concat: entity work.concat_c5804edea5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant4_op_net,
      in1 => mux_y_net_x0,
      in2 => addsub_s_net_x0,
      in3 => constant3_op_net,
      y => concat_y_net_x0
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net_x0
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net_x0
    );

  constant3: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_9f5572ba51
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant7: entity work.constant_c4c603edf2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net_x0
    );

  constant8: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net_x0
    );

  simulation_multiplexer: entity work.xlpassthrough
    generic map (
      din_width => 64,
      dout_width => 64
    )
    port map (
      din => bram_din_net_x0,
      dout => simulation_multiplexer_dout_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/BRAM IF 64b/Byte Sel"

entity byte_sel_entity_a0de3ec24a is
  port (
    b_sel: in std_logic_vector(2 downto 0); 
    x64b: in std_logic_vector(63 downto 0); 
    b: out std_logic_vector(7 downto 0)
  );
end byte_sel_entity_a0de3ec24a;

architecture structural of byte_sel_entity_a0de3ec24a is
  signal b0_y_net: std_logic_vector(7 downto 0);
  signal b1_y_net: std_logic_vector(7 downto 0);
  signal b2_y_net: std_logic_vector(7 downto 0);
  signal b3_y_net: std_logic_vector(7 downto 0);
  signal b4_y_net: std_logic_vector(7 downto 0);
  signal b5_y_net: std_logic_vector(7 downto 0);
  signal b6_y_net: std_logic_vector(7 downto 0);
  signal b7_y_net: std_logic_vector(7 downto 0);
  signal delay4_q_net_x0: std_logic_vector(2 downto 0);
  signal mux_y_net_x0: std_logic_vector(7 downto 0);
  signal simulation_multiplexer_dout_net_x1: std_logic_vector(63 downto 0);

begin
  delay4_q_net_x0 <= b_sel;
  simulation_multiplexer_dout_net_x1 <= x64b;
  b <= mux_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 32,
      new_msb => 39,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 47,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 48,
      new_msb => 55,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 56,
      new_msb => 63,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => simulation_multiplexer_dout_net_x1,
      y => b7_y_net
    );

  mux: entity work.mux_c762ea476a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b0_y_net,
      d1 => b1_y_net,
      d2 => b2_y_net,
      d3 => b3_y_net,
      d4 => b4_y_net,
      d5 => b5_y_net,
      d6 => b6_y_net,
      d7 => b7_y_net,
      sel => delay4_q_net_x0,
      y => mux_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/BRAM IF 64b"

entity bram_if_64b_entity_32e52dc467 is
  port (
    bram_din: in std_logic_vector(63 downto 0); 
    byte_addr: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    logical3: in std_logic; 
    regtx_pkt_buf_addr_offset: in std_logic_vector(7 downto 0); 
    tx_pkt_buf_sel: in std_logic_vector(3 downto 0); 
    bram_interface: out std_logic_vector(31 downto 0); 
    bram_interface_x0: out std_logic; 
    bram_interface_x1: out std_logic; 
    bram_interface_x2: out std_logic_vector(63 downto 0); 
    bram_interface_x3: out std_logic_vector(7 downto 0); 
    ram_byte: out std_logic_vector(7 downto 0)
  );
end bram_if_64b_entity_32e52dc467;

architecture structural of bram_if_64b_entity_32e52dc467 is
  signal addsub_s_net_x0: std_logic_vector(8 downto 0);
  signal bram_din_net_x1: std_logic_vector(63 downto 0);
  signal bytes_y_net_x2: std_logic_vector(11 downto 0);
  signal ce_1_sg_x38: std_logic;
  signal clk_1_sg_x38: std_logic;
  signal concat_y_net_x1: std_logic_vector(31 downto 0);
  signal constant1_op_net_x1: std_logic;
  signal constant2_op_net_x1: std_logic;
  signal constant7_op_net_x1: std_logic_vector(63 downto 0);
  signal constant8_op_net_x1: std_logic_vector(7 downto 0);
  signal delay4_q_net_x0: std_logic_vector(2 downto 0);
  signal logical3_y_net_x4: std_logic;
  signal mux5_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x2: std_logic_vector(3 downto 0);
  signal mux_y_net_x3: std_logic_vector(7 downto 0);
  signal n_msb_y_net: std_logic_vector(8 downto 0);
  signal register16_q_net_x0: std_logic_vector(7 downto 0);
  signal simulation_multiplexer_dout_net_x1: std_logic_vector(63 downto 0);
  signal x12_lsb_y_net_x0: std_logic_vector(11 downto 0);
  signal x3_lsb_y_net: std_logic_vector(2 downto 0);

begin
  bram_din_net_x1 <= bram_din;
  bytes_y_net_x2 <= byte_addr;
  ce_1_sg_x38 <= ce_1;
  clk_1_sg_x38 <= clk_1;
  logical3_y_net_x4 <= logical3;
  register16_q_net_x0 <= regtx_pkt_buf_addr_offset;
  mux_y_net_x2 <= tx_pkt_buf_sel;
  bram_interface <= concat_y_net_x1;
  bram_interface_x0 <= constant1_op_net_x1;
  bram_interface_x1 <= constant2_op_net_x1;
  bram_interface_x2 <= constant7_op_net_x1;
  bram_interface_x3 <= constant8_op_net_x1;
  ram_byte <= mux_y_net_x3;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 9,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 10,
      core_name0 => "addsb_11_0_73986f767e994888",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 10,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => register16_q_net_x0,
      b => n_msb_y_net,
      ce => ce_1_sg_x38,
      clk => clk_1_sg_x38,
      clr => '0',
      en => "1",
      s => addsub_s_net_x0
    );

  bram_addr_map_8b602ce2fb: entity work.bram_addr_map_entity_8b602ce2fb
    port map (
      ce_1 => ce_1_sg_x38,
      clk_1 => clk_1_sg_x38,
      tx_ind => x12_lsb_y_net_x0,
      tx_phy_mode_11n_ac => logical3_y_net_x4,
      mem_addr => mux5_y_net_x0
    );

  bram_interface_5cb2ccffdd: entity work.bram_interface_entity_5cb2ccffdd
    port map (
      bram_din => bram_din_net_x1,
      pkt_buf_index => mux_y_net_x2,
      x64b_word_addr => addsub_s_net_x0,
      concat_x0 => concat_y_net_x1,
      constant1_x0 => constant1_op_net_x1,
      constant2_x0 => constant2_op_net_x1,
      constant7_x0 => constant7_op_net_x1,
      constant8_x0 => constant8_op_net_x1,
      x64b_data => simulation_multiplexer_dout_net_x1
    );

  byte_sel_a0de3ec24a: entity work.byte_sel_entity_a0de3ec24a
    port map (
      b_sel => delay4_q_net_x0,
      x64b => simulation_multiplexer_dout_net_x1,
      b => mux_y_net_x3
    );

  delay4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 3
    )
    port map (
      ce => ce_1_sg_x38,
      clk => clk_1_sg_x38,
      d => x3_lsb_y_net,
      en => '1',
      rst => '1',
      q => delay4_q_net_x0
    );

  n_msb: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 11,
      x_width => 12,
      y_width => 9
    )
    port map (
      x => mux5_y_net_x0,
      y => n_msb_y_net
    );

  x12_lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 12,
      y_width => 12
    )
    port map (
      x => bytes_y_net_x2,
      y => x12_lsb_y_net_x0
    );

  x3_lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 12,
      y_width => 3
    )
    port map (
      x => mux5_y_net_x0,
      y => x3_lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/Bit Select"

entity bit_select_entity_4d6daa9b45 is
  port (
    b: in std_logic_vector(7 downto 0); 
    b_sel: in std_logic_vector(2 downto 0); 
    b_x0: out std_logic
  );
end bit_select_entity_4d6daa9b45;

architecture structural of bit_select_entity_4d6daa9b45 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b4_y_net: std_logic;
  signal b5_y_net: std_logic;
  signal b6_y_net: std_logic;
  signal b7_y_net: std_logic;
  signal delay5_q_net_x0: std_logic_vector(2 downto 0);
  signal mux1_y_net_x0: std_logic_vector(7 downto 0);
  signal mux_y_net_x0: std_logic;

begin
  mux1_y_net_x0 <= b;
  delay5_q_net_x0 <= b_sel;
  b_x0 <= mux_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux1_y_net_x0,
      y(0) => b7_y_net
    );

  mux: entity work.mux_b0082e75ff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b0_y_net,
      d1(0) => b1_y_net,
      d2(0) => b2_y_net,
      d3(0) => b3_y_net,
      d4(0) => b4_y_net,
      d5(0) => b5_y_net,
      d6(0) => b6_y_net,
      d7(0) => b7_y_net,
      sel => delay5_q_net_x0,
      y(0) => mux_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/Byte Src Sel"

entity byte_src_sel_entity_b4e477e100 is
  port (
    data_b: in std_logic_vector(7 downto 0); 
    fcs_b: in std_logic_vector(7 downto 0); 
    htsig: in std_logic_vector(7 downto 0); 
    sel_fcs: in std_logic; 
    sel_htsig: in std_logic; 
    sel_zero: in std_logic; 
    tx_byte: out std_logic_vector(7 downto 0)
  );
end byte_src_sel_entity_b4e477e100;

architecture structural of byte_src_sel_entity_b4e477e100 is
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant2_op_net: std_logic_vector(7 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay6_q_net_x0: std_logic;
  signal delay7_q_net_x0: std_logic;
  signal mux1_y_net_x1: std_logic_vector(7 downto 0);
  signal mux_y_net: std_logic_vector(7 downto 0);
  signal mux_y_net_x5: std_logic_vector(7 downto 0);
  signal mux_y_net_x6: std_logic_vector(7 downto 0);
  signal mux_y_net_x7: std_logic_vector(7 downto 0);

begin
  mux_y_net_x5 <= data_b;
  mux_y_net_x6 <= fcs_b;
  mux_y_net_x7 <= htsig;
  delay7_q_net_x0 <= sel_fcs;
  delay10_q_net_x0 <= sel_htsig;
  delay6_q_net_x0 <= sel_zero;
  tx_byte <= mux1_y_net_x1;

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay10_q_net_x0,
      in1(0) => delay7_q_net_x0,
      y => concat_y_net
    );

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  mux: entity work.mux_998e20a1ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux_y_net_x5,
      d1 => mux_y_net_x6,
      d2 => mux_y_net_x7,
      d3 => constant2_op_net,
      sel => concat_y_net,
      y => mux_y_net
    );

  mux1: entity work.mux_387191112d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux_y_net,
      d1 => constant1_op_net,
      sel(0) => delay6_q_net_x0,
      y => mux1_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/FCS Calc/Byte Sel"

entity byte_sel_entity_30fb4df82d is
  port (
    b_sel: in std_logic_vector(1 downto 0); 
    x32b: in std_logic_vector(31 downto 0); 
    b: out std_logic_vector(7 downto 0)
  );
end byte_sel_entity_30fb4df82d;

architecture structural of byte_sel_entity_30fb4df82d is
  signal addsub_s_net_x0: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(31 downto 0);
  signal b0_y_net: std_logic_vector(7 downto 0);
  signal b1_y_net: std_logic_vector(7 downto 0);
  signal b2_y_net: std_logic_vector(7 downto 0);
  signal b3_y_net: std_logic_vector(7 downto 0);
  signal mux_y_net_x7: std_logic_vector(7 downto 0);

begin
  addsub_s_net_x0 <= b_sel;
  assert_dout_net_x0 <= x32b;
  b <= mux_y_net_x7;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert_dout_net_x0,
      y => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert_dout_net_x0,
      y => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert_dout_net_x0,
      y => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert_dout_net_x0,
      y => b3_y_net
    );

  mux: entity work.mux_998e20a1ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b3_y_net,
      d1 => b2_y_net,
      d2 => b1_y_net,
      d3 => b0_y_net,
      sel => addsub_s_net_x0,
      y => mux_y_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/FCS Calc/CRC32 Calc/Endian Swap"

entity endian_swap_entity_da8729ff07 is
  port (
    b: in std_logic_vector(7 downto 0); 
    i: out std_logic_vector(7 downto 0)
  );
end endian_swap_entity_da8729ff07;

architecture structural of endian_swap_entity_da8729ff07 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b4_y_net: std_logic;
  signal b5_y_net: std_logic;
  signal b6_y_net: std_logic;
  signal b7_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal mux_y_net_x6: std_logic_vector(7 downto 0);

begin
  mux_y_net_x6 <= b;
  i <= concat_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x6,
      y(0) => b7_y_net
    );

  concat: entity work.concat_7673b9b993
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => b0_y_net,
      in1(0) => b1_y_net,
      in2(0) => b2_y_net,
      in3(0) => b3_y_net,
      in4(0) => b4_y_net,
      in5(0) => b5_y_net,
      in6(0) => b6_y_net,
      in7(0) => b7_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/FCS Calc/CRC32 Calc"

entity crc32_calc_entity_1f41b886a8 is
  port (
    byte: in std_logic_vector(7 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    tx_reset: in std_logic; 
    crc32: out std_logic_vector(31 downto 0)
  );
end crc32_calc_entity_1f41b886a8;

architecture structural of crc32_calc_entity_1f41b886a8 is
  signal assert1_dout_net: std_logic_vector(31 downto 0);
  signal assert_dout_net_x1: std_logic_vector(31 downto 0);
  signal b0_y_net_x1: std_logic_vector(7 downto 0);
  signal b1_y_net_x1: std_logic_vector(7 downto 0);
  signal b2_y_net_x1: std_logic_vector(7 downto 0);
  signal b3_y_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x39: std_logic;
  signal clk_1_sg_x39: std_logic;
  signal concat1_y_net: std_logic_vector(31 downto 0);
  signal concat_y_net: std_logic_vector(31 downto 0);
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concat_y_net_x2: std_logic_vector(7 downto 0);
  signal concat_y_net_x3: std_logic_vector(7 downto 0);
  signal concat_y_net_x4: std_logic_vector(7 downto 0);
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal crc_accum_q_net: std_logic_vector(31 downto 0);
  signal crc_remainders1_data_net: std_logic_vector(31 downto 0);
  signal inverter_op_net: std_logic_vector(31 downto 0);
  signal logical3_y_net: std_logic_vector(7 downto 0);
  signal logical3_y_net_x1: std_logic;
  signal logical4_y_net: std_logic_vector(31 downto 0);
  signal logical_y_net_x20: std_logic;
  signal mux_y_net_x7: std_logic_vector(7 downto 0);
  signal x24lsb_y_net: std_logic_vector(23 downto 0);
  signal x8msb_y_net: std_logic_vector(7 downto 0);

begin
  mux_y_net_x7 <= byte;
  ce_1_sg_x39 <= ce_1;
  clk_1_sg_x39 <= clk_1;
  logical3_y_net_x1 <= en;
  logical_y_net_x20 <= tx_reset;
  crc32 <= assert_dout_net_x1;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 32,
      dout_width => 32
    )
    port map (
      din => crc_accum_q_net,
      dout => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 32,
      dout_width => 32
    )
    port map (
      din => concat_y_net,
      dout => assert_dout_net_x1
    );

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b0_y_net_x1
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b1_y_net_x1
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b2_y_net_x1
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b3_y_net_x1
    );

  concat: entity work.concat_a1e126f11c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concat_y_net_x1,
      in1 => concat_y_net_x2,
      in2 => concat_y_net_x3,
      in3 => concat_y_net_x4,
      y => concat_y_net
    );

  concat1: entity work.concat_c048fbe4a5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => x24lsb_y_net,
      in1 => constant1_op_net,
      y => concat1_y_net
    );

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  crc_accum: entity work.xlregister
    generic map (
      d_width => 32,
      init_value => b"11111111111111111111111111111111"
    )
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      d => logical4_y_net,
      en(0) => logical3_y_net_x1,
      rst(0) => logical_y_net_x20,
      q => crc_accum_q_net
    );

  crc_remainders1: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 8,
      c_address_width => 8,
      c_width => 32,
      core_name0 => "dmg_72_134e91999cae8947",
      latency => 0
    )
    port map (
      addr => logical3_y_net,
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      en => "1",
      data => crc_remainders1_data_net
    );

  endian_swap1_096929c09a: entity work.endian_swap_entity_da8729ff07
    port map (
      b => b0_y_net_x1,
      i => concat_y_net_x1
    );

  endian_swap2_d4e79e08cf: entity work.endian_swap_entity_da8729ff07
    port map (
      b => b1_y_net_x1,
      i => concat_y_net_x2
    );

  endian_swap3_e1cec24f8a: entity work.endian_swap_entity_da8729ff07
    port map (
      b => b2_y_net_x1,
      i => concat_y_net_x3
    );

  endian_swap4_96f57d2581: entity work.endian_swap_entity_da8729ff07
    port map (
      b => b3_y_net_x1,
      i => concat_y_net_x4
    );

  endian_swap_da8729ff07: entity work.endian_swap_entity_da8729ff07
    port map (
      b => mux_y_net_x7,
      i => concat_y_net_x0
    );

  inverter: entity work.inverter_6a3d3dd4e5
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      ip => assert1_dout_net,
      op => inverter_op_net
    );

  logical3: entity work.logical_59f8d33339
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => x8msb_y_net,
      d1 => concat_y_net_x0,
      y => logical3_y_net
    );

  logical4: entity work.logical_b23aa74086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat1_y_net,
      d1 => crc_remainders1_data_net,
      y => logical4_y_net
    );

  x24lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 23,
      x_width => 32,
      y_width => 24
    )
    port map (
      x => assert1_dout_net,
      y => x24lsb_y_net
    );

  x8msb: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert1_dout_net,
      y => x8msb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/FCS Calc/posedge"

entity posedge_entity_73e633add7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end posedge_entity_73e633add7;

architecture structural of posedge_entity_73e633add7 is
  signal ce_1_sg_x40: std_logic;
  signal clk_1_sg_x40: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net_x0: std_logic;

begin
  ce_1_sg_x40 <= ce_1;
  clk_1_sg_x40 <= clk_1;
  logical2_y_net_x0 <= d;
  q <= logical1_y_net_x0;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      d(0) => logical2_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      clr => '0',
      ip(0) => delay_q_net,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical2_y_net_x0,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/FCS Calc"

entity fcs_calc_entity_6017d3d209 is
  port (
    byte: in std_logic_vector(7 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    byte_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fcs_sel: in std_logic; 
    tx_phy_mode_11ag: in std_logic; 
    tx_phy_mode_11n: in std_logic; 
    tx_reset: in std_logic; 
    crc_byte: out std_logic_vector(7 downto 0)
  );
end fcs_calc_entity_6017d3d209;

architecture structural of fcs_calc_entity_6017d3d209 is
  signal addsub_s_net_x0: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(31 downto 0);
  signal ce_1_sg_x41: std_logic;
  signal clk_1_sg_x41: std_logic;
  signal constant2_op_net: std_logic_vector(2 downto 0);
  signal constant3_op_net: std_logic_vector(3 downto 0);
  signal delay1_q_net_x0: std_logic_vector(11 downto 0);
  signal delay3_q_net_x0: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical5_y_net: std_logic;
  signal logical_y_net_x21: std_logic;
  signal mux_y_net_x10: std_logic_vector(7 downto 0);
  signal mux_y_net_x9: std_logic_vector(7 downto 0);
  signal register_q_net: std_logic_vector(1 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal slice1_y_net_x5: std_logic;
  signal slice_y_net_x2: std_logic;
  signal x2lsb_y_net: std_logic_vector(1 downto 0);

begin
  mux_y_net_x9 <= byte;
  delay1_q_net_x0 <= byte_ind;
  delay3_q_net_x0 <= byte_valid;
  ce_1_sg_x41 <= ce_1;
  clk_1_sg_x41 <= clk_1;
  logical2_y_net_x1 <= fcs_sel;
  slice_y_net_x2 <= tx_phy_mode_11ag;
  slice1_y_net_x5 <= tx_phy_mode_11n;
  logical_y_net_x21 <= tx_reset;
  crc_byte <= mux_y_net_x10;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_7925f33378f00f6a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => register_q_net,
      b => x2lsb_y_net,
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      clr => '0',
      en => "1",
      s => addsub_s_net_x0
    );

  byte_sel_30fb4df82d: entity work.byte_sel_entity_30fb4df82d
    port map (
      b_sel => addsub_s_net_x0,
      x32b => assert_dout_net_x1,
      b => mux_y_net_x10
    );

  constant2: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_c0ce4ae10c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  crc32_calc_1f41b886a8: entity work.crc32_calc_entity_1f41b886a8
    port map (
      byte => mux_y_net_x9,
      ce_1 => ce_1_sg_x41,
      clk_1 => clk_1_sg_x41,
      en => logical3_y_net_x1,
      tx_reset => logical_y_net_x21,
      crc32 => assert_dout_net_x1
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      clr => '0',
      ip(0) => logical2_y_net_x1,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical2_y_net,
      d1(0) => logical5_y_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice_y_net_x2,
      d1(0) => delay3_q_net_x0,
      d2(0) => relational2_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net,
      d1(0) => inverter_op_net,
      y(0) => logical3_y_net_x1
    );

  logical5: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x5,
      d1(0) => delay3_q_net_x0,
      d2(0) => relational1_op_net,
      y(0) => logical5_y_net
    );

  posedge_73e633add7: entity work.posedge_entity_73e633add7
    port map (
      ce_1 => ce_1_sg_x41,
      clk_1 => clk_1_sg_x41,
      d => logical2_y_net_x1,
      q => logical1_y_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 2,
      init_value => b"00"
    )
    port map (
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      d => x2lsb_y_net,
      en(0) => logical1_y_net_x0,
      rst(0) => logical_y_net_x21,
      q => register_q_net
    );

  relational1: entity work.relational_28e8664d0c
    port map (
      a => delay1_q_net_x0,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_ae4e737ca0
    port map (
      a => delay1_q_net_x0,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  x2lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => delay1_q_net_x0,
      y => x2lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/Packet Sections"

entity packet_sections_entity_1aaa2624ab is
  port (
    bit_sel: in std_logic_vector(2 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ofdm_tx_data_length: in std_logic_vector(15 downto 0); 
    tx_phy_mode_11n: in std_logic; 
    data_done: out std_logic; 
    sel_fcs: out std_logic; 
    sel_htsig: out std_logic; 
    sel_zero: out std_logic; 
    unscrambled: out std_logic
  );
end packet_sections_entity_1aaa2624ab;

architecture structural of packet_sections_entity_1aaa2624ab is
  signal addsub1_s_net: std_logic_vector(16 downto 0);
  signal addsub2_s_net: std_logic_vector(17 downto 0);
  signal addsub3_s_net: std_logic_vector(4 downto 0);
  signal bit_in_byte_y_net_x2: std_logic_vector(2 downto 0);
  signal bytes_y_net_x3: std_logic_vector(11 downto 0);
  signal ce_1_sg_x42: std_logic;
  signal clk_1_sg_x42: std_logic;
  signal constant1_op_net: std_logic_vector(2 downto 0);
  signal constant2_op_net: std_logic_vector(3 downto 0);
  signal constant3_op_net: std_logic_vector(2 downto 0);
  signal constant4_op_net: std_logic_vector(2 downto 0);
  signal constant5_op_net: std_logic_vector(2 downto 0);
  signal constant6_op_net: std_logic_vector(3 downto 0);
  signal constant7_op_net: std_logic_vector(3 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal mux8_y_net: std_logic_vector(3 downto 0);
  signal pad_x0: std_logic;
  signal register11_q_net_x0: std_logic_vector(15 downto 0);
  signal relational1_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational5_op_net: std_logic;
  signal relational6_op_net: std_logic;
  signal relational7_op_net: std_logic;
  signal sig_htsig: std_logic;
  signal slice1_y_net_x6: std_logic;
  signal tail: std_logic;

begin
  bit_in_byte_y_net_x2 <= bit_sel;
  bytes_y_net_x3 <= byte_ind;
  ce_1_sg_x42 <= ce_1;
  clk_1_sg_x42 <= clk_1;
  register11_q_net_x0 <= ofdm_tx_data_length;
  slice1_y_net_x6 <= tx_phy_mode_11n;
  data_done <= logical3_y_net_x0;
  sel_fcs <= logical2_y_net_x2;
  sel_htsig <= logical5_y_net_x0;
  sel_zero <= pad_x0;
  unscrambled <= logical1_y_net_x0;

  addsub1: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 5,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 16,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 17,
      core_name0 => "addsb_11_0_f66fe30ee2d0a6f0",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 17,
      latency => 1,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 17
    )
    port map (
      a => addsub3_s_net,
      b => register11_q_net_x0,
      ce => ce_1_sg_x42,
      clk => clk_1_sg_x42,
      clr => '0',
      en => "1",
      s => addsub1_s_net
    );

  addsub2: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 17,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 3,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 18,
      core_name0 => "addsb_11_0_6695c8a33176d3c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 18,
      latency => 1,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 0,
      s_width => 18
    )
    port map (
      a => addsub1_s_net,
      b => constant3_op_net,
      ce => ce_1_sg_x42,
      clk => clk_1_sg_x42,
      clr => '0',
      en => "1",
      s => addsub2_s_net
    );

  addsub3: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 4,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 3,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 5,
      core_name0 => "addsb_11_0_2fe7f24afe1bc972",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 5,
      latency => 1,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 5
    )
    port map (
      a => mux8_y_net,
      b => constant5_op_net,
      ce => ce_1_sg_x42,
      clk => clk_1_sg_x42,
      clr => '0',
      en => "1",
      s => addsub3_s_net
    );

  constant1: entity work.constant_0f59f02ba5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_a629aefb53
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_263f209841
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_1f5cc32f1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_a629aefb53
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  constant7: entity work.constant_8038205d89
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x42,
      clk => clk_1_sg_x42,
      clr => '0',
      ip(0) => pad_x0,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x42,
      clk => clk_1_sg_x42,
      clr => '0',
      ip(0) => relational6_op_net,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => sig_htsig,
      d1(0) => tail,
      y(0) => logical1_y_net_x0
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => relational1_op_net,
      y(0) => logical2_y_net_x2
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter1_op_net,
      d1(0) => relational5_op_net,
      y(0) => logical3_y_net_x0
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational6_op_net,
      d1(0) => relational5_op_net,
      y(0) => tail
    );

  logical5: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x6,
      d1(0) => relational3_op_net,
      d2(0) => relational7_op_net,
      y(0) => logical5_y_net_x0
    );

  mux8: entity work.mux_1e60cf48bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant1_op_net,
      d1 => constant2_op_net,
      sel(0) => slice1_y_net_x6,
      y => mux8_y_net
    );

  relational1: entity work.relational_82200c2969
    port map (
      a => bytes_y_net_x3,
      b => addsub2_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_31ab9f25e5
    port map (
      a => bytes_y_net_x3,
      b => mux8_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => sig_htsig
    );

  relational3: entity work.relational_31ab9f25e5
    port map (
      a => bytes_y_net_x3,
      b => constant6_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  relational4: entity work.relational_61c9d3f3fc
    port map (
      a => bytes_y_net_x3,
      b => addsub1_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_x0
    );

  relational5: entity work.relational_ab46f67027
    port map (
      a => bytes_y_net_x3,
      b => addsub1_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net
    );

  relational6: entity work.relational_6c709b1b0c
    port map (
      a => bit_in_byte_y_net_x2,
      b => constant4_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational6_op_net
    );

  relational7: entity work.relational_28e8664d0c
    port map (
      a => bytes_y_net_x3,
      b => constant7_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational7_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/CRC8 Calc/4LSB Calc"

entity x4lsb_calc_entity_a6845a4290 is
  port (
    crc_accum: in std_logic_vector(7 downto 0); 
    final_4lsb: out std_logic_vector(3 downto 0)
  );
end x4lsb_calc_entity_a6845a4290;

architecture structural of x4lsb_calc_entity_a6845a4290 is
  signal b_0_y_net: std_logic;
  signal b_1_y_net: std_logic;
  signal b_6_y_net: std_logic;
  signal b_7_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(3 downto 0);
  signal crc_accum_q_net_x0: std_logic_vector(7 downto 0);
  signal logical1_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;

begin
  crc_accum_q_net_x0 <= crc_accum;
  final_4lsb <= concat_y_net_x0;

  b_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => crc_accum_q_net_x0,
      y(0) => b_0_y_net
    );

  b_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => crc_accum_q_net_x0,
      y(0) => b_1_y_net
    );

  b_6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => crc_accum_q_net_x0,
      y(0) => b_6_y_net
    );

  b_7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => crc_accum_q_net_x0,
      y(0) => b_7_y_net
    );

  concat: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => logical3_y_net,
      in1(0) => logical4_y_net,
      in2(0) => logical1_y_net,
      in3(0) => b_6_y_net,
      y => concat_y_net_x0
    );

  logical1: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b_6_y_net,
      d1(0) => b_7_y_net,
      y(0) => logical1_y_net
    );

  logical3: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b_1_y_net,
      d1(0) => b_7_y_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b_0_y_net,
      d1(0) => logical1_y_net,
      y(0) => logical4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/CRC8 Calc"

entity crc8_calc_entity_023caf907a is
  port (
    byte_ind: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_byte: in std_logic_vector(7 downto 0); 
    data_valid: in std_logic; 
    reset: in std_logic; 
    crc8: out std_logic_vector(7 downto 0)
  );
end crc8_calc_entity_023caf907a;

architecture structural of crc8_calc_entity_023caf907a is
  signal assert1_dout_net: std_logic_vector(7 downto 0);
  signal b_5_2_y_net: std_logic_vector(3 downto 0);
  signal ce_1_sg_x43: std_logic;
  signal clk_1_sg_x43: std_logic;
  signal concat3_y_net: std_logic_vector(7 downto 0);
  signal concat_y_net_x0: std_logic_vector(3 downto 0);
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal constant3_op_net: std_logic_vector(3 downto 0);
  signal constant4_op_net: std_logic_vector(3 downto 0);
  signal crc8_lookup_data_net: std_logic_vector(7 downto 0);
  signal crc_accum_q_net_x0: std_logic_vector(7 downto 0);
  signal delay1_q_net_x1: std_logic_vector(11 downto 0);
  signal delay3_q_net_x1: std_logic;
  signal inverter_op_net_x0: std_logic_vector(7 downto 0);
  signal logical1_y_net: std_logic;
  signal logical3_y_net: std_logic_vector(7 downto 0);
  signal logical_y_net_x22: std_logic;
  signal mux_y_net_x11: std_logic_vector(7 downto 0);
  signal relational3_op_net: std_logic;
  signal relational4_op_net: std_logic;

begin
  delay1_q_net_x1 <= byte_ind;
  ce_1_sg_x43 <= ce_1;
  clk_1_sg_x43 <= clk_1;
  mux_y_net_x11 <= data_byte;
  delay3_q_net_x1 <= data_valid;
  logical_y_net_x22 <= reset;
  crc8 <= inverter_op_net_x0;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 8,
      dout_width => 8
    )
    port map (
      din => crc_accum_q_net_x0,
      dout => assert1_dout_net
    );

  b_5_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 5,
      x_width => 8,
      y_width => 4
    )
    port map (
      x => assert1_dout_net,
      y => b_5_2_y_net
    );

  concat3: entity work.concat_1a070f1f35
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => b_5_2_y_net,
      in1 => concat_y_net_x0,
      y => concat3_y_net
    );

  constant3: entity work.constant_8038205d89
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_bfd5ba0f50
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  crc8_lookup: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 8,
      c_address_width => 8,
      c_width => 8,
      core_name0 => "dmg_72_06262d82a068201e",
      latency => 0
    )
    port map (
      addr => logical3_y_net,
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      en => "1",
      data => crc8_lookup_data_net
    );

  crc_accum: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"11111111"
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => crc8_lookup_data_net,
      en(0) => logical1_y_net,
      rst(0) => logical_y_net_x22,
      q => crc_accum_q_net_x0
    );

  endian_swap_8c480d3f51: entity work.endian_swap_entity_da8729ff07
    port map (
      b => mux_y_net_x11,
      i => concat_y_net_x1
    );

  inverter: entity work.inverter_4a6def08e4
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip => concat3_y_net,
      op => inverter_op_net_x0
    );

  logical1: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x1,
      d1(0) => relational3_op_net,
      d2(0) => relational4_op_net,
      y(0) => logical1_y_net
    );

  logical3: entity work.logical_59f8d33339
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => assert1_dout_net,
      d1 => concat_y_net_x1,
      y => logical3_y_net
    );

  relational3: entity work.relational_28e8664d0c
    port map (
      a => delay1_q_net_x1,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  relational4: entity work.relational_b218b04ee6
    port map (
      a => delay1_q_net_x1,
      b => constant4_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  x4lsb_calc_a6845a4290: entity work.x4lsb_calc_entity_a6845a4290
    port map (
      crc_accum => crc_accum_q_net_x0,
      final_4lsb => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/Format"

entity format_entity_0ad24997d8 is
  port (
    crc: in std_logic_vector(7 downto 0); 
    htsig_4: out std_logic_vector(7 downto 0); 
    htsig_5: out std_logic_vector(7 downto 0)
  );
end format_entity_0ad24997d8;

architecture structural of format_entity_0ad24997d8 is
  signal b_1_0_y_net: std_logic_vector(1 downto 0);
  signal b_7_2_y_net: std_logic_vector(5 downto 0);
  signal concat1_y_net_x0: std_logic_vector(7 downto 0);
  signal concat2_y_net_x0: std_logic_vector(7 downto 0);
  signal concat_y_net_x2: std_logic_vector(7 downto 0);
  signal concat_y_net_x3: std_logic_vector(7 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal inverter_op_net_x1: std_logic_vector(7 downto 0);

begin
  inverter_op_net_x1 <= crc;
  htsig_4 <= concat_y_net_x2;
  htsig_5 <= concat_y_net_x3;

  b_1_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => inverter_op_net_x1,
      y => b_1_0_y_net
    );

  b_7_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 7,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => inverter_op_net_x1,
      y => b_7_2_y_net
    );

  concat1: entity work.concat_dc245eb1d2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => b_1_0_y_net,
      in1 => constant2_op_net,
      y => concat1_y_net_x0
    );

  concat2: entity work.concat_dc245eb1d2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant1_op_net,
      in1 => b_7_2_y_net,
      y => concat2_y_net_x0
    );

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_7ea0f2fff7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  endian_swap1_6bd84470ea: entity work.endian_swap_entity_da8729ff07
    port map (
      b => concat2_y_net_x0,
      i => concat_y_net_x2
    );

  endian_swap2_de497d11a4: entity work.endian_swap_entity_da8729ff07
    port map (
      b => concat1_y_net_x0,
      i => concat_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/HT Length"

entity ht_length_entity_07f41e4db8 is
  port (
    b4: in std_logic_vector(7 downto 0); 
    b5: in std_logic_vector(7 downto 0); 
    length: out std_logic_vector(15 downto 0)
  );
end ht_length_entity_07f41e4db8;

architecture structural of ht_length_entity_07f41e4db8 is
  signal concat1_y_net_x0: std_logic_vector(15 downto 0);
  signal dout1_q_net_x0: std_logic_vector(7 downto 0);
  signal dout2_q_net_x0: std_logic_vector(7 downto 0);

begin
  dout1_q_net_x0 <= b4;
  dout2_q_net_x0 <= b5;
  length <= concat1_y_net_x0;

  concat1: entity work.concat_8e53793314
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => dout2_q_net_x0,
      in1 => dout1_q_net_x0,
      y => concat1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/HT-SIG Flags"

entity ht_sig_flags_entity_129b03e671 is
  port (
    b3: in std_logic_vector(7 downto 0); 
    b6: in std_logic_vector(7 downto 0); 
    b7: in std_logic_vector(7 downto 0); 
    unsupported: out std_logic
  );
end ht_sig_flags_entity_129b03e671;

architecture structural of ht_sig_flags_entity_129b03e671 is
  signal b_1_0_y_net: std_logic_vector(1 downto 0);
  signal b_5_4_y_net: std_logic_vector(1 downto 0);
  signal b_6_y_net: std_logic;
  signal b_7_y_net: std_logic;
  signal b_7_y_net_x0: std_logic;
  signal constant1_op_net: std_logic;
  signal constant_op_net: std_logic;
  signal dout3_q_net_x0: std_logic_vector(7 downto 0);
  signal dout4_q_net_x0: std_logic_vector(7 downto 0);
  signal dout_q_net_x0: std_logic_vector(7 downto 0);
  signal logical_y_net_x0: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  dout_q_net_x0 <= b3;
  dout3_q_net_x0 <= b6;
  dout4_q_net_x0 <= b7;
  unsupported <= logical_y_net_x0;

  b_1_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => dout4_q_net_x0,
      y => b_1_0_y_net
    );

  b_5_4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 5,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => dout3_q_net_x0,
      y => b_5_4_y_net
    );

  b_6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout3_q_net_x0,
      y(0) => b_6_y_net
    );

  b_7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x0,
      y(0) => b_7_y_net
    );

  b_7_x0: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout3_q_net_x0,
      y(0) => b_7_y_net_x0
    );

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant_x0: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  logical: entity work.logical_0ee569a826
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b_7_y_net,
      d1(0) => b_6_y_net,
      d2(0) => b_7_y_net_x0,
      d3(0) => relational1_op_net,
      d4(0) => relational_op_net,
      y(0) => logical_y_net_x0
    );

  relational: entity work.relational_2a3f3bef9d
    port map (
      a => b_1_0_y_net,
      b(0) => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_2a3f3bef9d
    port map (
      a => b_5_4_y_net,
      b(0) => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode/MCS Decode"

entity mcs_decode_entity_39140b24b4 is
  port (
    b3: in std_logic_vector(7 downto 0); 
    b6: in std_logic_vector(7 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    code_rate: out std_logic_vector(1 downto 0); 
    mcs_valid: out std_logic; 
    mod_sel: out std_logic_vector(1 downto 0); 
    n_dbps: out std_logic_vector(9 downto 0); 
    unsupported: out std_logic
  );
end mcs_decode_entity_39140b24b4;

architecture structural of mcs_decode_entity_39140b24b4 is
  signal b_0_y_net: std_logic;
  signal b_26_17_y_net: std_logic_vector(9 downto 0);
  signal b_4_3_y_net: std_logic_vector(1 downto 0);
  signal b_6_5_y_net: std_logic_vector(1 downto 0);
  signal b_7_y_net: std_logic;
  signal ce_1_sg_x44: std_logic;
  signal clk_1_sg_x44: std_logic;
  signal concat_y_net: std_logic_vector(5 downto 0);
  signal constant17_op_net: std_logic_vector(2 downto 0);
  signal constant18_op_net: std_logic_vector(6 downto 0);
  signal convert_dout_net: std_logic;
  signal dout3_q_net_x1: std_logic_vector(7 downto 0);
  signal dout_q_net_x1: std_logic_vector(7 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal relational_op_net: std_logic;
  signal rom_data_net: std_logic_vector(31 downto 0);
  signal x5lsb_y_net: std_logic_vector(4 downto 0);
  signal x7lsb_y_net: std_logic_vector(6 downto 0);

begin
  dout_q_net_x1 <= b3;
  dout3_q_net_x1 <= b6;
  ce_1_sg_x44 <= ce_1;
  clk_1_sg_x44 <= clk_1;
  code_rate <= b_6_5_y_net;
  mcs_valid <= relational1_op_net_x0;
  mod_sel <= b_4_3_y_net;
  n_dbps <= b_26_17_y_net;
  unsupported <= logical1_y_net_x0;

  b_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => rom_data_net,
      y(0) => b_0_y_net
    );

  b_26_17: entity work.xlslice
    generic map (
      new_lsb => 17,
      new_msb => 26,
      x_width => 32,
      y_width => 10
    )
    port map (
      x => rom_data_net,
      y => b_26_17_y_net
    );

  b_4_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 32,
      y_width => 2
    )
    port map (
      x => rom_data_net,
      y => b_4_3_y_net
    );

  b_6_5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 32,
      y_width => 2
    )
    port map (
      x => rom_data_net,
      y => b_6_5_y_net
    );

  b_7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout3_q_net_x1,
      y(0) => b_7_y_net
    );

  concat: entity work.concat_ac785d9b37
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => b_7_y_net,
      in1 => x5lsb_y_net,
      y => concat_y_net
    );

  constant17: entity work.constant_1d6ad1c713
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant17_op_net
    );

  constant18: entity work.constant_1a631d900c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant18_op_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      clr => '0',
      din(0) => b_0_y_net,
      en => "1",
      dout(0) => convert_dout_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert_dout_net,
      d1(0) => relational_op_net,
      y(0) => logical1_y_net_x0
    );

  relational: entity work.relational_c5ffb0182e
    port map (
      a => x7lsb_y_net,
      b => constant17_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_27dbff5dcf
    port map (
      a => x7lsb_y_net,
      b => constant18_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  rom: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 6,
      c_width => 32,
      core_name0 => "bmg_72_d44417b0abe027bf",
      latency => 1
    )
    port map (
      addr => concat_y_net,
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      en => "1",
      rst => "0",
      data => rom_data_net
    );

  x5lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 8,
      y_width => 5
    )
    port map (
      x => dout_q_net_x1,
      y => x5lsb_y_net
    );

  x7lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 6,
      x_width => 8,
      y_width => 7
    )
    port map (
      x => dout_q_net_x1,
      y => x7lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/HT-SIG Decode"

entity ht_sig_decode_entity_aae4465e4a is
  port (
    byte: in std_logic_vector(7 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    byte_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    rst: in std_logic; 
    code_rate: out std_logic_vector(1 downto 0); 
    ht_sig_bytes: out std_logic_vector(7 downto 0); 
    ht_sig_invalid: out std_logic; 
    ht_sig_valid: out std_logic; 
    length: out std_logic_vector(15 downto 0); 
    mod_sel: out std_logic_vector(1 downto 0); 
    n_dbps: out std_logic_vector(9 downto 0); 
    unsupported: out std_logic
  );
end ht_sig_decode_entity_aae4465e4a;

architecture structural of ht_sig_decode_entity_aae4465e4a is
  signal b_26_17_y_net_x0: std_logic_vector(9 downto 0);
  signal b_4_3_y_net_x0: std_logic_vector(1 downto 0);
  signal b_6_5_y_net_x0: std_logic_vector(1 downto 0);
  signal ce_1_sg_x45: std_logic;
  signal clk_1_sg_x45: std_logic;
  signal concat1_y_net_x1: std_logic_vector(15 downto 0);
  signal concat2_y_net: std_logic_vector(1 downto 0);
  signal concat_y_net_x2: std_logic_vector(7 downto 0);
  signal concat_y_net_x3: std_logic_vector(7 downto 0);
  signal constant1_op_net: std_logic_vector(2 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic_vector(2 downto 0);
  signal constant4_op_net: std_logic_vector(3 downto 0);
  signal constant5_op_net: std_logic_vector(2 downto 0);
  signal constant_op_net: std_logic_vector(2 downto 0);
  signal delay1_q_net: std_logic;
  signal delay1_q_net_x2: std_logic_vector(11 downto 0);
  signal delay3_q_net_x2: std_logic;
  signal delay_q_net: std_logic;
  signal dout1_q_net_x0: std_logic_vector(7 downto 0);
  signal dout2_q_net_x0: std_logic_vector(7 downto 0);
  signal dout3_q_net_x1: std_logic_vector(7 downto 0);
  signal dout4_q_net_x0: std_logic_vector(7 downto 0);
  signal dout_q_net_x1: std_logic_vector(7 downto 0);
  signal inverter4_op_net: std_logic;
  signal inverter_op_net_x1: std_logic_vector(7 downto 0);
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;
  signal logical5_y_net: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal logical9_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x23: std_logic;
  signal mux_y_net_x12: std_logic_vector(7 downto 0);
  signal mux_y_net_x8: std_logic_vector(7 downto 0);
  signal relational1_op_net: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational4_op_net: std_logic;
  signal relational5_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  mux_y_net_x12 <= byte;
  delay1_q_net_x2 <= byte_ind;
  delay3_q_net_x2 <= byte_valid;
  ce_1_sg_x45 <= ce_1;
  clk_1_sg_x45 <= clk_1;
  logical_y_net_x23 <= rst;
  code_rate <= b_6_5_y_net_x0;
  ht_sig_bytes <= mux_y_net_x8;
  ht_sig_invalid <= logical6_y_net_x0;
  ht_sig_valid <= logical8_y_net_x0;
  length <= concat1_y_net_x1;
  mod_sel <= b_4_3_y_net_x0;
  n_dbps <= b_26_17_y_net_x0;
  unsupported <= logical9_y_net_x0;

  concat2: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => relational3_op_net,
      in1(0) => relational4_op_net,
      y => concat2_y_net
    );

  constant1: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_1d6ad1c713
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_145086465d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_263f209841
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant_x0: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  crc8_calc_023caf907a: entity work.crc8_calc_entity_023caf907a
    port map (
      byte_ind => delay1_q_net_x2,
      ce_1 => ce_1_sg_x45,
      clk_1 => clk_1_sg_x45,
      data_byte => mux_y_net_x12,
      data_valid => delay3_q_net_x2,
      reset => logical_y_net_x23,
      crc8 => inverter_op_net_x1
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d(0) => logical3_y_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d(0) => delay_q_net,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  dout: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d => mux_y_net_x12,
      en(0) => logical2_y_net,
      rst(0) => logical_y_net_x23,
      q => dout_q_net_x1
    );

  dout1: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"01100100"
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d => mux_y_net_x12,
      en(0) => logical1_y_net,
      rst(0) => logical_y_net_x23,
      q => dout1_q_net_x0
    );

  dout2: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d => mux_y_net_x12,
      en(0) => logical_y_net,
      rst(0) => logical_y_net_x23,
      q => dout2_q_net_x0
    );

  dout3: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000011"
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d => mux_y_net_x12,
      en(0) => logical5_y_net,
      rst(0) => logical_y_net_x23,
      q => dout3_q_net_x1
    );

  dout4: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"11100000"
    )
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      d => mux_y_net_x12,
      en(0) => logical4_y_net,
      rst(0) => logical_y_net_x23,
      q => dout4_q_net_x0
    );

  format_0ad24997d8: entity work.format_entity_0ad24997d8
    port map (
      crc => inverter_op_net_x1,
      htsig_4 => concat_y_net_x2,
      htsig_5 => concat_y_net_x3
    );

  ht_length_07f41e4db8: entity work.ht_length_entity_07f41e4db8
    port map (
      b4 => dout1_q_net_x0,
      b5 => dout2_q_net_x0,
      length => concat1_y_net_x1
    );

  ht_sig_flags_129b03e671: entity work.ht_sig_flags_entity_129b03e671
    port map (
      b3 => dout_q_net_x1,
      b6 => dout3_q_net_x1,
      b7 => dout4_q_net_x0,
      unsupported => logical_y_net_x0
    );

  inverter4: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x45,
      clk => clk_1_sg_x45,
      clr => '0',
      ip(0) => relational1_op_net_x0,
      op(0) => inverter4_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational_op_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational4_op_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational3_op_net,
      y(0) => logical4_y_net
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x2,
      d1(0) => relational5_op_net,
      y(0) => logical5_y_net
    );

  logical6: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter4_op_net,
      d1(0) => delay1_q_net,
      y(0) => logical6_y_net_x0
    );

  logical8: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x0,
      d1(0) => delay1_q_net,
      y(0) => logical8_y_net_x0
    );

  logical9: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x0,
      d1(0) => logical_y_net_x0,
      y(0) => logical9_y_net_x0
    );

  mcs_decode_39140b24b4: entity work.mcs_decode_entity_39140b24b4
    port map (
      b3 => dout_q_net_x1,
      b6 => dout3_q_net_x1,
      ce_1 => ce_1_sg_x45,
      clk_1 => clk_1_sg_x45,
      code_rate => b_6_5_y_net_x0,
      mcs_valid => relational1_op_net_x0,
      mod_sel => b_4_3_y_net_x0,
      n_dbps => b_26_17_y_net_x0,
      unsupported => logical1_y_net_x0
    );

  mux: entity work.mux_f1cd62c228
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux_y_net_x12,
      d1 => concat_y_net_x3,
      d2 => concat_y_net_x2,
      sel => concat2_y_net,
      y => mux_y_net_x8
    );

  relational: entity work.relational_09ceb5d9bd
    port map (
      a => delay1_q_net_x2,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_09ceb5d9bd
    port map (
      a => delay1_q_net_x2,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_ae8b814968
    port map (
      a => delay1_q_net_x2,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_09ceb5d9bd
    port map (
      a => delay1_q_net_x2,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  relational4: entity work.relational_5321bc1192
    port map (
      a => delay1_q_net_x2,
      b => constant4_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  relational5: entity work.relational_09ceb5d9bd
    port map (
      a => delay1_q_net_x2,
      b => constant5_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode/LENGTH"

entity length_entity_8cda74b311 is
  port (
    b0: in std_logic_vector(7 downto 0); 
    b1: in std_logic_vector(7 downto 0); 
    b2: in std_logic_vector(7 downto 0); 
    length: out std_logic_vector(11 downto 0)
  );
end length_entity_8cda74b311;

architecture structural of length_entity_8cda74b311 is
  signal concat_y_net_x0: std_logic_vector(11 downto 0);
  signal dout1_q_net_x0: std_logic_vector(7 downto 0);
  signal dout2_q_net_x0: std_logic_vector(7 downto 0);
  signal dout_q_net_x0: std_logic_vector(7 downto 0);
  signal x1lsb_y_net: std_logic;
  signal x3msb_y_net: std_logic_vector(2 downto 0);

begin
  dout_q_net_x0 <= b0;
  dout1_q_net_x0 <= b1;
  dout2_q_net_x0 <= b2;
  length <= concat_y_net_x0;

  concat: entity work.concat_1d9bdbb01e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => x1lsb_y_net,
      in1 => dout1_q_net_x0,
      in2 => x3msb_y_net,
      y => concat_y_net_x0
    );

  x1lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout2_q_net_x0,
      y(0) => x1lsb_y_net
    );

  x3msb: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 7,
      x_width => 8,
      y_width => 3
    )
    port map (
      x => dout_q_net_x0,
      y => x3msb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode/RATE Decode"

entity rate_decode_entity_3797b32f88 is
  port (
    b0: in std_logic_vector(7 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    code_rate: out std_logic_vector(1 downto 0); 
    mod_sel: out std_logic_vector(1 downto 0); 
    n_dbps: out std_logic_vector(9 downto 0); 
    rate_valid: out std_logic
  );
end rate_decode_entity_3797b32f88;

architecture structural of rate_decode_entity_3797b32f88 is
  signal b_26_17_y_net: std_logic_vector(9 downto 0);
  signal b_4_3_y_net: std_logic_vector(1 downto 0);
  signal b_6_5_y_net: std_logic_vector(1 downto 0);
  signal ce_1_sg_x47: std_logic;
  signal clk_1_sg_x47: std_logic;
  signal constant17_op_net: std_logic_vector(2 downto 0);
  signal constant18_op_net: std_logic_vector(2 downto 0);
  signal constant19_op_net: std_logic_vector(2 downto 0);
  signal constant20_op_net: std_logic_vector(2 downto 0);
  signal constant21_op_net: std_logic_vector(2 downto 0);
  signal constant22_op_net: std_logic_vector(2 downto 0);
  signal constant23_op_net: std_logic_vector(2 downto 0);
  signal constant24_op_net: std_logic_vector(2 downto 0);
  signal dout_q_net_x1: std_logic_vector(7 downto 0);
  signal msb_y_net_x0: std_logic;
  signal mux3_y_net: std_logic_vector(2 downto 0);
  signal rom_data_net: std_logic_vector(31 downto 0);
  signal x3lsb_y_net: std_logic_vector(2 downto 0);
  signal x4lsb_y_net: std_logic_vector(3 downto 0);

begin
  dout_q_net_x1 <= b0;
  ce_1_sg_x47 <= ce_1;
  clk_1_sg_x47 <= clk_1;
  code_rate <= b_6_5_y_net;
  mod_sel <= b_4_3_y_net;
  n_dbps <= b_26_17_y_net;
  rate_valid <= msb_y_net_x0;

  b_26_17: entity work.xlslice
    generic map (
      new_lsb => 17,
      new_msb => 26,
      x_width => 32,
      y_width => 10
    )
    port map (
      x => rom_data_net,
      y => b_26_17_y_net
    );

  b_4_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 32,
      y_width => 2
    )
    port map (
      x => rom_data_net,
      y => b_4_3_y_net
    );

  b_6_5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 32,
      y_width => 2
    )
    port map (
      x => rom_data_net,
      y => b_6_5_y_net
    );

  constant17: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant17_op_net
    );

  constant18: entity work.constant_a1c496ea88
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant18_op_net
    );

  constant19: entity work.constant_1f5cc32f1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant19_op_net
    );

  constant20: entity work.constant_0f59f02ba5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant20_op_net
    );

  constant21: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant21_op_net
    );

  constant22: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant22_op_net
    );

  constant23: entity work.constant_263f209841
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant23_op_net
    );

  constant24: entity work.constant_1d6ad1c713
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant24_op_net
    );

  msb: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => x4lsb_y_net,
      y(0) => msb_y_net_x0
    );

  mux3: entity work.mux_8a8a6c93e0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant23_op_net,
      d1 => constant21_op_net,
      d2 => constant19_op_net,
      d3 => constant17_op_net,
      d4 => constant24_op_net,
      d5 => constant22_op_net,
      d6 => constant20_op_net,
      d7 => constant18_op_net,
      sel => x3lsb_y_net,
      y => mux3_y_net
    );

  rom: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 3,
      c_width => 32,
      core_name0 => "bmg_72_8bdf24f02e925a98",
      latency => 1
    )
    port map (
      addr => mux3_y_net,
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      en => "1",
      rst => "0",
      data => rom_data_net
    );

  x3lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 4,
      y_width => 3
    )
    port map (
      x => x4lsb_y_net,
      y => x3lsb_y_net
    );

  x4lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 8,
      y_width => 4
    )
    port map (
      x => dout_q_net_x1,
      y => x4lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode/Tail & Parity Check/2b XOR"

entity x2b_xor_entity_a508f1e574 is
  port (
    a: in std_logic_vector(1 downto 0); 
    b: out std_logic
  );
end x2b_xor_entity_a508f1e574;

architecture structural of x2b_xor_entity_a508f1e574 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal x2lsb_y_net_x0: std_logic_vector(1 downto 0);

begin
  x2lsb_y_net_x0 <= a;
  b <= logical_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => x2lsb_y_net_x0,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => x2lsb_y_net_x0,
      y(0) => b1_y_net
    );

  logical: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b0_y_net,
      d1(0) => b1_y_net,
      y(0) => logical_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode/Tail & Parity Check/8b XOR 1"

entity x8b_xor_1_entity_ea024c6d09 is
  port (
    a: in std_logic_vector(7 downto 0); 
    b: out std_logic
  );
end x8b_xor_1_entity_ea024c6d09;

architecture structural of x8b_xor_1_entity_ea024c6d09 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b4_y_net: std_logic;
  signal b5_y_net: std_logic;
  signal b6_y_net: std_logic;
  signal b7_y_net: std_logic;
  signal dout_q_net_x2: std_logic_vector(7 downto 0);
  signal logical_y_net_x0: std_logic;

begin
  dout_q_net_x2 <= a;
  b <= logical_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => dout_q_net_x2,
      y(0) => b7_y_net
    );

  logical: entity work.logical_9ac2bdb119
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b0_y_net,
      d1(0) => b1_y_net,
      d2(0) => b2_y_net,
      d3(0) => b3_y_net,
      d4(0) => b4_y_net,
      d5(0) => b5_y_net,
      d6(0) => b6_y_net,
      d7(0) => b7_y_net,
      y(0) => logical_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode/Tail & Parity Check"

entity \tail___parity_check_entity_b17def6b42\ is
  port (
    b0: in std_logic_vector(7 downto 0); 
    b1: in std_logic_vector(7 downto 0); 
    b2: in std_logic_vector(7 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    invalid: out std_logic
  );
end \tail___parity_check_entity_b17def6b42\;

architecture structural of \tail___parity_check_entity_b17def6b42\ is
  signal ce_1_sg_x48: std_logic;
  signal clk_1_sg_x48: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal convert1_dout_net: std_logic;
  signal dout1_q_net_x2: std_logic_vector(7 downto 0);
  signal dout2_q_net_x1: std_logic_vector(7 downto 0);
  signal dout_q_net_x3: std_logic_vector(7 downto 0);
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x1: std_logic;
  signal logical_y_net_x2: std_logic;
  signal relational1_op_net: std_logic;
  signal x2lsb_y_net_x0: std_logic_vector(1 downto 0);
  signal x6msb_y_net: std_logic_vector(5 downto 0);

begin
  dout_q_net_x3 <= b0;
  dout1_q_net_x2 <= b1;
  dout2_q_net_x1 <= b2;
  ce_1_sg_x48 <= ce_1;
  clk_1_sg_x48 <= clk_1;
  invalid <= logical5_y_net_x0;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      clr => '0',
      din(0) => logical_y_net,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical: entity work.logical_604045dd09
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x1,
      d1(0) => logical_y_net_x2,
      d2(0) => logical_y_net_x0,
      y(0) => logical_y_net
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => relational1_op_net,
      y(0) => logical5_y_net_x0
    );

  relational1: entity work.relational_c49d820dc8
    port map (
      a => x6msb_y_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  x2b_xor_a508f1e574: entity work.x2b_xor_entity_a508f1e574
    port map (
      a => x2lsb_y_net_x0,
      b => logical_y_net_x0
    );

  x2lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => dout2_q_net_x1,
      y => x2lsb_y_net_x0
    );

  x6msb: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 7,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => dout2_q_net_x1,
      y => x6msb_y_net
    );

  x8b_xor_1_ea024c6d09: entity work.x8b_xor_1_entity_ea024c6d09
    port map (
      a => dout_q_net_x3,
      b => logical_y_net_x1
    );

  x8b_xor_2_960b7f64c7: entity work.x8b_xor_1_entity_ea024c6d09
    port map (
      a => dout1_q_net_x2,
      b => logical_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode/SIGNAL Decode"

entity signal_decode_entity_b2c8f51d1d is
  port (
    byte: in std_logic_vector(7 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    byte_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    rst: in std_logic; 
    code_rate: out std_logic_vector(1 downto 0); 
    length: out std_logic_vector(11 downto 0); 
    mod_sel: out std_logic_vector(1 downto 0); 
    n_dbps: out std_logic_vector(9 downto 0); 
    signal_invalid: out std_logic
  );
end signal_decode_entity_b2c8f51d1d;

architecture structural of signal_decode_entity_b2c8f51d1d is
  signal b_26_17_y_net_x0: std_logic_vector(9 downto 0);
  signal b_4_3_y_net_x0: std_logic_vector(1 downto 0);
  signal b_6_5_y_net_x0: std_logic_vector(1 downto 0);
  signal ce_1_sg_x49: std_logic;
  signal clk_1_sg_x49: std_logic;
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x3: std_logic_vector(11 downto 0);
  signal delay3_q_net_x3: std_logic;
  signal delay_q_net: std_logic;
  signal dout1_q_net_x2: std_logic_vector(7 downto 0);
  signal dout2_q_net_x1: std_logic_vector(7 downto 0);
  signal dout_q_net_x3: std_logic_vector(7 downto 0);
  signal inverter3_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical5_y_net: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x25: std_logic;
  signal msb_y_net_x0: std_logic;
  signal mux_y_net_x13: std_logic_vector(7 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  mux_y_net_x13 <= byte;
  delay1_q_net_x3 <= byte_ind;
  delay3_q_net_x3 <= byte_valid;
  ce_1_sg_x49 <= ce_1;
  clk_1_sg_x49 <= clk_1;
  logical_y_net_x25 <= rst;
  code_rate <= b_6_5_y_net_x0;
  length <= concat_y_net_x1;
  mod_sel <= b_4_3_y_net_x0;
  n_dbps <= b_26_17_y_net_x0;
  signal_invalid <= logical3_y_net_x0;

  constant1: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant_x0: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x49,
      clk => clk_1_sg_x49,
      d(0) => logical_y_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  dout: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"01101011"
    )
    port map (
      ce => ce_1_sg_x49,
      clk => clk_1_sg_x49,
      d => mux_y_net_x13,
      en(0) => logical2_y_net,
      rst(0) => logical_y_net_x25,
      q => dout_q_net_x3
    );

  dout1: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000111"
    )
    port map (
      ce => ce_1_sg_x49,
      clk => clk_1_sg_x49,
      d => mux_y_net_x13,
      en(0) => logical1_y_net,
      rst(0) => logical_y_net_x25,
      q => dout1_q_net_x2
    );

  dout2: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x49,
      clk => clk_1_sg_x49,
      d => mux_y_net_x13,
      en(0) => logical_y_net,
      rst(0) => logical_y_net_x25,
      q => dout2_q_net_x1
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x49,
      clk => clk_1_sg_x49,
      clr => '0',
      ip(0) => msb_y_net_x0,
      op(0) => inverter3_op_net
    );

  length_8cda74b311: entity work.length_entity_8cda74b311
    port map (
      b0 => dout_q_net_x3,
      b1 => dout1_q_net_x2,
      b2 => dout2_q_net_x1,
      length => concat_y_net_x1
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x3,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x3,
      d1(0) => relational_op_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay3_q_net_x3,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net,
      d1(0) => logical5_y_net,
      y(0) => logical3_y_net_x0
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter3_op_net,
      d1(0) => logical5_y_net_x0,
      y(0) => logical5_y_net
    );

  rate_decode_3797b32f88: entity work.rate_decode_entity_3797b32f88
    port map (
      b0 => dout_q_net_x3,
      ce_1 => ce_1_sg_x49,
      clk_1 => clk_1_sg_x49,
      code_rate => b_6_5_y_net_x0,
      mod_sel => b_4_3_y_net_x0,
      n_dbps => b_26_17_y_net_x0,
      rate_valid => msb_y_net_x0
    );

  relational: entity work.relational_ae8b814968
    port map (
      a => delay1_q_net_x3,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_ae8b814968
    port map (
      a => delay1_q_net_x3,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_ae8b814968
    port map (
      a => delay1_q_net_x3,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  tail_parity_check_b17def6b42: entity work.\tail___parity_check_entity_b17def6b42\
    port map (
      b0 => dout_q_net_x3,
      b1 => dout1_q_net_x2,
      b2 => dout2_q_net_x1,
      ce_1 => ce_1_sg_x49,
      clk_1 => clk_1_sg_x49,
      invalid => logical5_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/SIGNAL & HT-SIG Decode"

entity \signal___ht_sig_decode_entity_18bbc6a95e\ is
  port (
    byte: in std_logic_vector(7 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    tx_phy_mode_11n: in std_logic; 
    tx_reset: in std_logic; 
    valid: in std_logic; 
    ht_sig_bytes: out std_logic_vector(7 downto 0); 
    ofdm_tx_data_code_rate: out std_logic_vector(1 downto 0); 
    ofdm_tx_data_length: out std_logic_vector(15 downto 0); 
    ofdm_tx_data_mod_sel: out std_logic_vector(1 downto 0); 
    ofdm_tx_data_n_dbps: out std_logic_vector(9 downto 0); 
    reset_phy: out std_logic
  );
end \signal___ht_sig_decode_entity_18bbc6a95e\;

architecture structural of \signal___ht_sig_decode_entity_18bbc6a95e\ is
  signal b_26_17_y_net_x0: std_logic_vector(9 downto 0);
  signal b_26_17_y_net_x1: std_logic_vector(9 downto 0);
  signal b_4_3_y_net_x0: std_logic_vector(1 downto 0);
  signal b_4_3_y_net_x1: std_logic_vector(1 downto 0);
  signal b_6_5_y_net_x0: std_logic_vector(1 downto 0);
  signal b_6_5_y_net_x1: std_logic_vector(1 downto 0);
  signal ce_1_sg_x50: std_logic;
  signal clk_1_sg_x50: std_logic;
  signal concat1_y_net_x1: std_logic_vector(15 downto 0);
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal delay1_q_net_x4: std_logic_vector(11 downto 0);
  signal delay3_q_net_x4: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical4_y_net_x0: std_logic;
  signal logical5_y_net: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal logical9_y_net_x0: std_logic;
  signal logical_y_net_x26: std_logic;
  signal mux2_y_net: std_logic_vector(9 downto 0);
  signal mux3_y_net: std_logic_vector(15 downto 0);
  signal mux7_y_net: std_logic_vector(1 downto 0);
  signal mux8_y_net: std_logic_vector(1 downto 0);
  signal mux_y_net_x14: std_logic_vector(7 downto 0);
  signal mux_y_net_x9: std_logic_vector(7 downto 0);
  signal register11_q_net_x1: std_logic_vector(15 downto 0);
  signal register1_q_net_x2: std_logic_vector(9 downto 0);
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x2: std_logic_vector(1 downto 0);
  signal register3_q_net_x0: std_logic_vector(1 downto 0);
  signal slice1_y_net_x7: std_logic;

begin
  mux_y_net_x14 <= byte;
  delay1_q_net_x4 <= byte_ind;
  ce_1_sg_x50 <= ce_1;
  clk_1_sg_x50 <= clk_1;
  slice1_y_net_x7 <= tx_phy_mode_11n;
  logical_y_net_x26 <= tx_reset;
  delay3_q_net_x4 <= valid;
  ht_sig_bytes <= mux_y_net_x9;
  ofdm_tx_data_code_rate <= register3_q_net_x0;
  ofdm_tx_data_length <= register11_q_net_x1;
  ofdm_tx_data_mod_sel <= register2_q_net_x2;
  ofdm_tx_data_n_dbps <= register1_q_net_x2;
  reset_phy <= logical4_y_net_x0;

  ht_sig_decode_aae4465e4a: entity work.ht_sig_decode_entity_aae4465e4a
    port map (
      byte => mux_y_net_x14,
      byte_ind => delay1_q_net_x4,
      byte_valid => delay3_q_net_x4,
      ce_1 => ce_1_sg_x50,
      clk_1 => clk_1_sg_x50,
      rst => logical_y_net_x26,
      code_rate => b_6_5_y_net_x0,
      ht_sig_bytes => mux_y_net_x9,
      ht_sig_invalid => logical6_y_net_x0,
      ht_sig_valid => logical8_y_net_x0,
      length => concat1_y_net_x1,
      mod_sel => b_4_3_y_net_x0,
      n_dbps => b_26_17_y_net_x0,
      unsupported => logical9_y_net_x0
    );

  logical1: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x7,
      d1(0) => logical8_y_net_x0,
      d2(0) => logical9_y_net_x0,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical8_y_net_x0,
      d1(0) => slice1_y_net_x7,
      y(0) => logical2_y_net_x0
    );

  logical4: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical3_y_net_x0,
      d1(0) => logical1_y_net,
      d2(0) => logical5_y_net,
      y(0) => logical4_y_net_x0
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x7,
      d1(0) => logical6_y_net_x0,
      y(0) => logical5_y_net
    );

  mux2: entity work.mux_eb88ab7682
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b_26_17_y_net_x1,
      d1 => b_26_17_y_net_x0,
      sel(0) => register2_q_net_x1,
      y => mux2_y_net
    );

  mux3: entity work.mux_a585e6d5ba
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat_y_net_x1,
      d1 => concat1_y_net_x1,
      sel(0) => register2_q_net_x1,
      y => mux3_y_net
    );

  mux7: entity work.mux_2a63ac73aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b_6_5_y_net_x1,
      d1 => b_6_5_y_net_x0,
      sel(0) => register2_q_net_x1,
      y => mux7_y_net
    );

  mux8: entity work.mux_2a63ac73aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b_4_3_y_net_x1,
      d1 => b_4_3_y_net_x0,
      sel(0) => register2_q_net_x1,
      y => mux8_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 10,
      init_value => b"0000000000"
    )
    port map (
      ce => ce_1_sg_x50,
      clk => clk_1_sg_x50,
      d => mux2_y_net,
      en => "1",
      rst => "0",
      q => register1_q_net_x2
    );

  register11: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x50,
      clk => clk_1_sg_x50,
      d => mux3_y_net,
      en => "1",
      rst => "0",
      q => register11_q_net_x1
    );

  register2: entity work.xlregister
    generic map (
      d_width => 2,
      init_value => b"00"
    )
    port map (
      ce => ce_1_sg_x50,
      clk => clk_1_sg_x50,
      d => mux8_y_net,
      en => "1",
      rst => "0",
      q => register2_q_net_x2
    );

  register3: entity work.xlregister
    generic map (
      d_width => 2,
      init_value => b"00"
    )
    port map (
      ce => ce_1_sg_x50,
      clk => clk_1_sg_x50,
      d => mux7_y_net,
      en => "1",
      rst => "0",
      q => register3_q_net_x0
    );

  s_r_latch1_3ced5309b4: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x50,
      clk_1 => clk_1_sg_x50,
      r => logical_y_net_x26,
      s => logical2_y_net_x0,
      q => register2_q_net_x1
    );

  signal_decode_b2c8f51d1d: entity work.signal_decode_entity_b2c8f51d1d
    port map (
      byte => mux_y_net_x14,
      byte_ind => delay1_q_net_x4,
      byte_valid => delay3_q_net_x4,
      ce_1 => ce_1_sg_x50,
      clk_1 => clk_1_sg_x50,
      rst => logical_y_net_x26,
      code_rate => b_6_5_y_net_x1,
      length => concat_y_net_x1,
      mod_sel => b_4_3_y_net_x1,
      n_dbps => b_26_17_y_net_x1,
      signal_invalid => logical3_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/Scrambling/Scrambling LFSR"

entity scrambling_lfsr_entity_2d0e0f870d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    regtx_reset_scrambling_lfsr_perpkt: in std_logic; 
    tx_reset: in std_logic; 
    q: out std_logic
  );
end scrambling_lfsr_entity_2d0e0f870d;

architecture structural of scrambling_lfsr_entity_2d0e0f870d is
  signal assert1_dout_net: std_logic;
  signal assert_dout_net: std_logic;
  signal ce_1_sg_x51: std_logic;
  signal clk_1_sg_x51: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x27: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register6_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x51 <= ce_1;
  clk_1_sg_x51 <= clk_1;
  logical2_y_net_x0 <= en;
  register2_q_net_x1 <= regtx_reset_scrambling_lfsr_perpkt;
  logical_y_net_x27 <= tx_reset;
  q <= convert2_dout_net_x0;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register3_q_net,
      dout(0) => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register6_q_net,
      dout(0) => assert_dout_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      clr => '0',
      din(0) => logical1_y_net,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      clr => '0',
      din(0) => logical2_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      clr => '0',
      din(0) => logical_y_net,
      en => "1",
      dout(0) => convert2_dout_net_x0
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => assert_dout_net,
      d1(0) => assert1_dout_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x27,
      d1(0) => register2_q_net_x1,
      y(0) => logical1_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register1_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register2_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register3_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register4_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => register5_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register6_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x51,
      clk => clk_1_sg_x51,
      d(0) => logical_y_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/Scrambling"

entity scrambling_entity_cb9b9374d7 is
  port (
    bit: in std_logic; 
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    logical_x0: in std_logic; 
    register2: in std_logic; 
    unscrambled: in std_logic; 
    tx_bit: out std_logic
  );
end scrambling_entity_cb9b9374d7;

architecture structural of scrambling_entity_cb9b9374d7 is
  signal ce_1_sg_x52: std_logic;
  signal clk_1_sg_x52: std_logic;
  signal convert2_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal delay2_q_net_x2: std_logic;
  signal delay4_q_net_x0: std_logic;
  signal inverter1_op_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net: std_logic;
  signal logical_y_net_x1: std_logic;
  signal logical_y_net_x28: std_logic;
  signal mux_y_net_x1: std_logic;
  signal register2_q_net_x2: std_logic;

begin
  mux_y_net_x1 <= bit;
  delay2_q_net_x2 <= bit_valid;
  ce_1_sg_x52 <= ce_1;
  clk_1_sg_x52 <= clk_1;
  logical_y_net_x28 <= logical_x0;
  register2_q_net_x2 <= register2;
  delay4_q_net_x0 <= unscrambled;
  tx_bit <= logical_y_net_x1;

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x52,
      clk => clk_1_sg_x52,
      clr => '0',
      din(0) => inverter1_op_net,
      en => "1",
      dout(0) => convert2_dout_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x52,
      clk => clk_1_sg_x52,
      clr => '0',
      ip(0) => delay4_q_net_x0,
      op(0) => inverter1_op_net
    );

  logical: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical3_y_net,
      d1(0) => mux_y_net_x1,
      y(0) => logical_y_net_x1
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net_x2,
      d1(0) => inverter1_op_net,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert2_dout_net_x0,
      d1(0) => convert2_dout_net,
      y(0) => logical3_y_net
    );

  scrambling_lfsr_2d0e0f870d: entity work.scrambling_lfsr_entity_2d0e0f870d
    port map (
      ce_1 => ce_1_sg_x52,
      clk_1 => clk_1_sg_x52,
      en => logical2_y_net_x0,
      regtx_reset_scrambling_lfsr_perpkt => register2_q_net_x2,
      tx_reset => logical_y_net_x28,
      q => convert2_dout_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data/negedge"

entity negedge_entity_1004c64c9c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end negedge_entity_1004c64c9c;

architecture structural of negedge_entity_1004c64c9c is
  signal ce_1_sg_x53: std_logic;
  signal clk_1_sg_x53: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical4_y_net_x3: std_logic;

begin
  ce_1_sg_x53 <= ce_1;
  clk_1_sg_x53 <= clk_1;
  logical4_y_net_x3 <= d;
  q <= logical1_y_net_x1;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d(0) => logical4_y_net_x3,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      clr => '0',
      ip(0) => logical4_y_net_x3,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => delay_q_net,
      y(0) => logical1_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Pkt Data"

entity pkt_data_entity_6db78f9ff0 is
  port (
    bit_sel: in std_logic_vector(2 downto 0); 
    bit_sel_valid: in std_logic; 
    bram_din: in std_logic_vector(63 downto 0); 
    byte_ind: in std_logic_vector(11 downto 0); 
    byte_ind_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    logical: in std_logic; 
    logical3: in std_logic; 
    mux: in std_logic_vector(3 downto 0); 
    register16: in std_logic_vector(7 downto 0); 
    register2: in std_logic; 
    slice: in std_logic; 
    slice1: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    bram_if_64b: out std_logic_vector(31 downto 0); 
    bram_if_64b_x0: out std_logic; 
    bram_if_64b_x1: out std_logic; 
    bram_if_64b_x2: out std_logic_vector(63 downto 0); 
    bram_if_64b_x3: out std_logic_vector(7 downto 0); 
    data_done: out std_logic; 
    signal_ht_sig_decode: out std_logic_vector(9 downto 0); 
    signal_ht_sig_decode_x0: out std_logic_vector(1 downto 0); 
    signal_ht_sig_decode_x1: out std_logic_vector(1 downto 0); 
    sym_cfg_x0: out std_logic_vector(17 downto 0); 
    tx_bit: out std_logic; 
    tx_bit_tlast: out std_logic; 
    tx_bit_tvalid: out std_logic; 
    tx_sig_decode_error: out std_logic
  );
end pkt_data_entity_6db78f9ff0;

architecture structural of pkt_data_entity_6db78f9ff0 is
  signal bit_in_byte_y_net_x3: std_logic_vector(2 downto 0);
  signal bram_din_net_x2: std_logic_vector(63 downto 0);
  signal bytes_y_net_x4: std_logic_vector(11 downto 0);
  signal ce_1_sg_x54: std_logic;
  signal clk_1_sg_x54: std_logic;
  signal concat_y_net_x2: std_logic_vector(31 downto 0);
  signal concat_y_net_x6: std_logic_vector(17 downto 0);
  signal constant1_op_net_x2: std_logic;
  signal constant2_op_net_x2: std_logic;
  signal constant7_op_net_x2: std_logic_vector(63 downto 0);
  signal constant8_op_net_x2: std_logic_vector(7 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x4: std_logic_vector(11 downto 0);
  signal delay2_q_net_x3: std_logic;
  signal delay3_q_net_x4: std_logic;
  signal delay4_q_net_x0: std_logic;
  signal delay5_q_net_x0: std_logic_vector(2 downto 0);
  signal delay6_q_net_x0: std_logic;
  signal delay7_q_net_x0: std_logic;
  signal delay8_q_net_x1: std_logic_vector(17 downto 0);
  signal delay9_q_net_x2: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical3_y_net_x5: std_logic;
  signal logical4_y_net_x4: std_logic;
  signal logical4_y_net_x5: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical5_y_net_x2: std_logic;
  signal logical_y_net_x2: std_logic;
  signal logical_y_net_x29: std_logic;
  signal mux1_y_net_x1: std_logic_vector(7 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x10: std_logic_vector(7 downto 0);
  signal mux_y_net_x11: std_logic_vector(3 downto 0);
  signal mux_y_net_x14: std_logic_vector(7 downto 0);
  signal mux_y_net_x9: std_logic_vector(7 downto 0);
  signal pad_x0: std_logic;
  signal register11_q_net_x1: std_logic_vector(15 downto 0);
  signal register16_q_net_x1: std_logic_vector(7 downto 0);
  signal register1_q_net_x3: std_logic_vector(9 downto 0);
  signal register2_q_net_x4: std_logic;
  signal register2_q_net_x5: std_logic_vector(1 downto 0);
  signal register3_q_net_x1: std_logic_vector(1 downto 0);
  signal slice1_y_net_x8: std_logic;
  signal slice_y_net_x3: std_logic;

begin
  bit_in_byte_y_net_x3 <= bit_sel;
  logical4_y_net_x4 <= bit_sel_valid;
  bram_din_net_x2 <= bram_din;
  bytes_y_net_x4 <= byte_ind;
  logical5_y_net_x2 <= byte_ind_valid;
  ce_1_sg_x54 <= ce_1;
  clk_1_sg_x54 <= clk_1;
  logical_y_net_x29 <= logical;
  logical3_y_net_x5 <= logical3;
  mux_y_net_x11 <= mux;
  register16_q_net_x1 <= register16;
  register2_q_net_x4 <= register2;
  slice_y_net_x3 <= slice;
  slice1_y_net_x8 <= slice1;
  concat_y_net_x6 <= sym_cfg;
  bram_if_64b <= concat_y_net_x2;
  bram_if_64b_x0 <= constant1_op_net_x2;
  bram_if_64b_x1 <= constant2_op_net_x2;
  bram_if_64b_x2 <= constant7_op_net_x2;
  bram_if_64b_x3 <= constant8_op_net_x2;
  data_done <= delay9_q_net_x2;
  signal_ht_sig_decode <= register1_q_net_x3;
  signal_ht_sig_decode_x0 <= register2_q_net_x5;
  signal_ht_sig_decode_x1 <= register3_q_net_x1;
  sym_cfg_x0 <= delay8_q_net_x1;
  tx_bit <= logical_y_net_x2;
  tx_bit_tlast <= logical1_y_net_x2;
  tx_bit_tvalid <= delay2_q_net_x3;
  tx_sig_decode_error <= logical4_y_net_x5;

  bit_select_4d6daa9b45: entity work.bit_select_entity_4d6daa9b45
    port map (
      b => mux1_y_net_x1,
      b_sel => delay5_q_net_x0,
      b_x0 => mux_y_net_x1
    );

  bram_if_64b_32e52dc467: entity work.bram_if_64b_entity_32e52dc467
    port map (
      bram_din => bram_din_net_x2,
      byte_addr => bytes_y_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      logical3 => logical3_y_net_x5,
      regtx_pkt_buf_addr_offset => register16_q_net_x1,
      tx_pkt_buf_sel => mux_y_net_x11,
      bram_interface => concat_y_net_x2,
      bram_interface_x0 => constant1_op_net_x2,
      bram_interface_x1 => constant2_op_net_x2,
      bram_interface_x2 => constant7_op_net_x2,
      bram_interface_x3 => constant8_op_net_x2,
      ram_byte => mux_y_net_x14
    );

  byte_src_sel_b4e477e100: entity work.byte_src_sel_entity_b4e477e100
    port map (
      data_b => mux_y_net_x14,
      fcs_b => mux_y_net_x10,
      htsig => mux_y_net_x9,
      sel_fcs => delay7_q_net_x0,
      sel_htsig => delay10_q_net_x0,
      sel_zero => delay6_q_net_x0,
      tx_byte => mux1_y_net_x1
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d => bytes_y_net_x4,
      en => '1',
      rst => '1',
      q => delay1_q_net_x4
    );

  delay10: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical5_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay10_q_net_x0
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical4_y_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x3
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical5_y_net_x2,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x4
    );

  delay4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay4_q_net_x0
    );

  delay5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 3
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d => bit_in_byte_y_net_x3,
      en => '1',
      rst => '1',
      q => delay5_q_net_x0
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => pad_x0,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net_x0
    );

  delay7: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical2_y_net_x2,
      en => '1',
      rst => '1',
      q(0) => delay7_q_net_x0
    );

  delay8: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d => concat_y_net_x6,
      en => '1',
      rst => '1',
      q => delay8_q_net_x1
    );

  delay9: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      d(0) => logical3_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay9_q_net_x2
    );

  fcs_calc_6017d3d209: entity work.fcs_calc_entity_6017d3d209
    port map (
      byte => mux_y_net_x14,
      byte_ind => delay1_q_net_x4,
      byte_valid => delay3_q_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      fcs_sel => logical2_y_net_x2,
      tx_phy_mode_11ag => slice_y_net_x3,
      tx_phy_mode_11n => slice1_y_net_x8,
      tx_reset => logical_y_net_x29,
      crc_byte => mux_y_net_x10
    );

  negedge_1004c64c9c: entity work.negedge_entity_1004c64c9c
    port map (
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      d => logical4_y_net_x4,
      q => logical1_y_net_x2
    );

  packet_sections_1aaa2624ab: entity work.packet_sections_entity_1aaa2624ab
    port map (
      bit_sel => bit_in_byte_y_net_x3,
      byte_ind => bytes_y_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      ofdm_tx_data_length => register11_q_net_x1,
      tx_phy_mode_11n => slice1_y_net_x8,
      data_done => logical3_y_net_x0,
      sel_fcs => logical2_y_net_x2,
      sel_htsig => logical5_y_net_x0,
      sel_zero => pad_x0,
      unscrambled => logical1_y_net_x0
    );

  scrambling_cb9b9374d7: entity work.scrambling_entity_cb9b9374d7
    port map (
      bit => mux_y_net_x1,
      bit_valid => delay2_q_net_x3,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      logical_x0 => logical_y_net_x29,
      register2 => register2_q_net_x4,
      unscrambled => delay4_q_net_x0,
      tx_bit => logical_y_net_x2
    );

  signal_ht_sig_decode_18bbc6a95e: entity work.\signal___ht_sig_decode_entity_18bbc6a95e\
    port map (
      byte => mux_y_net_x14,
      byte_ind => delay1_q_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      tx_phy_mode_11n => slice1_y_net_x8,
      tx_reset => logical_y_net_x29,
      valid => delay3_q_net_x4,
      ht_sig_bytes => mux_y_net_x9,
      ofdm_tx_data_code_rate => register3_q_net_x1,
      ofdm_tx_data_length => register11_q_net_x1,
      ofdm_tx_data_mod_sel => register2_q_net_x5,
      ofdm_tx_data_n_dbps => register1_q_net_x3,
      reset_phy => logical4_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleave RAM"

entity interleave_ram_entity_42ac73a366 is
  port (
    bit_a: in std_logic; 
    bit_addr_a: in std_logic_vector(8 downto 0); 
    bit_addr_b: in std_logic_vector(8 downto 0); 
    bit_b: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    rd_addr: in std_logic_vector(5 downto 0); 
    rd_mem_sel: in std_logic; 
    wr_a: in std_logic; 
    wr_b: in std_logic; 
    wr_mem_sel: in std_logic; 
    sc_bits: out std_logic_vector(7 downto 0)
  );
end interleave_ram_entity_42ac73a366;

architecture structural of interleave_ram_entity_42ac73a366 is
  component interleaver_ram
    port (
      addra: in std_logic_vector(8 downto 0); 
      addrb: in std_logic_vector(8 downto 0); 
      ce: in std_logic; 
      clk: in std_logic; 
      dina: in std_logic_vector(0 downto 0); 
      dinb: in std_logic_vector(0 downto 0); 
      wea: in std_logic_vector(0 downto 0); 
      web: in std_logic_vector(0 downto 0); 
      douta: out std_logic_vector(7 downto 0); 
      doutb: out std_logic_vector(7 downto 0)
    );
  end component;
  signal assert1_dout_net: std_logic_vector(8 downto 0);
  signal assert_dout_net: std_logic_vector(8 downto 0);
  signal ce_1_sg_x55: std_logic;
  signal clk_1_sg_x55: std_logic;
  signal concat_y_net: std_logic_vector(8 downto 0);
  signal constant_op_net: std_logic_vector(2 downto 0);
  signal delay1_q_net_x1: std_logic;
  signal delay1_q_net_x2: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay2_q_net_x2: std_logic;
  signal interleaver_ram_0_douta_net: std_logic_vector(7 downto 0);
  signal interleaver_ram_0_doutb_net: std_logic_vector(7 downto 0);
  signal interleaver_ram_1_douta_net: std_logic_vector(7 downto 0);
  signal interleaver_ram_1_doutb_net: std_logic_vector(7 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter_op_net_x0: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;
  signal map_rom_douta_net_x0: std_logic_vector(8 downto 0);
  signal map_rom_doutb_net_x0: std_logic_vector(8 downto 0);
  signal mux1_y_net_x6: std_logic_vector(7 downto 0);
  signal mux2_y_net: std_logic_vector(8 downto 0);
  signal mux3_y_net: std_logic_vector(8 downto 0);
  signal register2_q_net_x0: std_logic;
  signal slice_y_net_x3: std_logic_vector(5 downto 0);

begin
  delay1_q_net_x1 <= bit_a;
  map_rom_douta_net_x0 <= bit_addr_a;
  map_rom_doutb_net_x0 <= bit_addr_b;
  delay2_q_net_x1 <= bit_b;
  ce_1_sg_x55 <= ce_1;
  clk_1_sg_x55 <= clk_1;
  slice_y_net_x3 <= rd_addr;
  register2_q_net_x0 <= rd_mem_sel;
  delay1_q_net_x2 <= wr_a;
  delay2_q_net_x2 <= wr_b;
  inverter_op_net_x0 <= wr_mem_sel;
  sc_bits <= mux1_y_net_x6;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 9,
      dout_width => 9
    )
    port map (
      din => mux3_y_net,
      dout => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 9,
      dout_width => 9
    )
    port map (
      din => mux2_y_net,
      dout => assert_dout_net
    );

  concat: entity work.concat_13241d6573
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => slice_y_net_x3,
      in1 => constant_op_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  interleaver_ram_0: interleaver_ram
    port map (
      addra => assert_dout_net,
      addrb => map_rom_doutb_net_x0,
      ce => ce_1_sg_x55,
      clk => clk_1_sg_x55,
      dina(0) => delay1_q_net_x1,
      dinb(0) => delay2_q_net_x1,
      wea(0) => logical3_y_net,
      web(0) => logical1_y_net,
      douta => interleaver_ram_0_douta_net,
      doutb => interleaver_ram_0_doutb_net
    );

  interleaver_ram_1: interleaver_ram
    port map (
      addra => assert1_dout_net,
      addrb => map_rom_doutb_net_x0,
      ce => ce_1_sg_x55,
      clk => clk_1_sg_x55,
      dina(0) => delay1_q_net_x1,
      dinb(0) => delay2_q_net_x1,
      wea(0) => logical4_y_net,
      web(0) => logical2_y_net,
      douta => interleaver_ram_1_douta_net,
      doutb => interleaver_ram_1_doutb_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x55,
      clk => clk_1_sg_x55,
      clr => '0',
      ip(0) => inverter_op_net_x0,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter1_op_net,
      d1(0) => delay2_q_net_x2,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net_x0,
      d1(0) => delay2_q_net_x2,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay1_q_net_x2,
      d1(0) => inverter1_op_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay1_q_net_x2,
      d1(0) => inverter_op_net_x0,
      y(0) => logical4_y_net
    );

  mux1: entity work.mux_387191112d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => interleaver_ram_0_douta_net,
      d1 => interleaver_ram_1_douta_net,
      sel(0) => register2_q_net_x0,
      y => mux1_y_net_x6
    );

  mux2: entity work.mux_791081a00e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat_y_net,
      d1 => map_rom_douta_net_x0,
      sel(0) => logical3_y_net,
      y => mux2_y_net
    );

  mux3: entity work.mux_791081a00e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat_y_net,
      d1 => map_rom_douta_net_x0,
      sel(0) => logical4_y_net,
      y => mux3_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Bit Index Calc"

entity bit_index_calc_entity_ec83e953ec is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    inc: in std_logic_vector(1 downto 0); 
    rst: in std_logic; 
    ind_a: out std_logic_vector(8 downto 0); 
    ind_b: out std_logic_vector(8 downto 0)
  );
end bit_index_calc_entity_ec83e953ec;

architecture structural of bit_index_calc_entity_ec83e953ec is
  signal accumulator_q_net_x0: std_logic_vector(8 downto 0);
  signal addsub_s_net_x0: std_logic_vector(8 downto 0);
  signal ce_1_sg_x56: std_logic;
  signal clk_1_sg_x56: std_logic;
  signal constant2_op_net: std_logic;
  signal delay3_q_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal mux4_y_net_x0: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x56 <= ce_1;
  clk_1_sg_x56 <= clk_1;
  delay3_q_net_x1 <= en;
  mux4_y_net_x0 <= inc;
  logical2_y_net_x0 <= rst;
  ind_a <= accumulator_q_net_x0;
  ind_b <= addsub_s_net_x0;

  accumulator: entity work.accum_3520344abf
    port map (
      b => mux4_y_net_x0,
      ce => ce_1_sg_x56,
      clk => clk_1_sg_x56,
      clr => '0',
      en(0) => delay3_q_net_x1,
      rst(0) => logical2_y_net_x0,
      q => accumulator_q_net_x0
    );

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 9,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 1,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 10,
      core_name0 => "addsb_11_0_73986f767e994888",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 10,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => accumulator_q_net_x0,
      b(0) => constant2_op_net,
      ce => ce_1_sg_x56,
      clk => clk_1_sg_x56,
      clr => '0',
      en => "1",
      s => addsub_s_net_x0
    );

  constant2: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Interleave Mapping"

entity interleave_mapping_entity_48a573e6d3 is
  port (
    base_rate_sym: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ind_a: in std_logic_vector(8 downto 0); 
    ind_b: in std_logic_vector(8 downto 0); 
    ofdm_tx_data_mod_sel: in std_logic_vector(1 downto 0); 
    tx_phy_mode_11n: in std_logic; 
    addr_a: out std_logic_vector(8 downto 0); 
    addr_b: out std_logic_vector(8 downto 0)
  );
end interleave_mapping_entity_48a573e6d3;

architecture structural of interleave_mapping_entity_48a573e6d3 is
  signal accumulator_q_net_x1: std_logic_vector(8 downto 0);
  signal addsub_s_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x57: std_logic;
  signal clk_1_sg_x57: std_logic;
  signal concat1_y_net: std_logic_vector(1 downto 0);
  signal concat2_y_net: std_logic_vector(11 downto 0);
  signal concat3_y_net: std_logic_vector(11 downto 0);
  signal constant8_op_net: std_logic_vector(8 downto 0);
  signal constant9_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net: std_logic_vector(1 downto 0);
  signal logical_y_net: std_logic;
  signal map_rom_douta_net_x1: std_logic_vector(8 downto 0);
  signal map_rom_doutb_net_x1: std_logic_vector(8 downto 0);
  signal mcode_load_base_rate_net_x0: std_logic;
  signal register2_q_net_x6: std_logic_vector(1 downto 0);
  signal slice1_y_net_x9: std_logic;

begin
  mcode_load_base_rate_net_x0 <= base_rate_sym;
  ce_1_sg_x57 <= ce_1;
  clk_1_sg_x57 <= clk_1;
  accumulator_q_net_x1 <= ind_a;
  addsub_s_net_x1 <= ind_b;
  register2_q_net_x6 <= ofdm_tx_data_mod_sel;
  slice1_y_net_x9 <= tx_phy_mode_11n;
  addr_a <= map_rom_douta_net_x1;
  addr_b <= map_rom_doutb_net_x1;

  concat1: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => inverter_op_net,
      in1(0) => inverter_op_net,
      y => concat1_y_net
    );

  concat2: entity work.concat_2d0bbe9efa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => logical_y_net,
      in1 => logical1_y_net,
      in2 => accumulator_q_net_x1,
      y => concat2_y_net
    );

  concat3: entity work.concat_2d0bbe9efa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => logical_y_net,
      in1 => logical1_y_net,
      in2 => addsub_s_net_x1,
      y => concat3_y_net
    );

  constant8: entity work.constant_fd85eb7067
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net
    );

  constant9: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant9_op_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      clr => '0',
      ip(0) => mcode_load_base_rate_net_x0,
      op(0) => inverter_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x9,
      d1(0) => inverter_op_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_33c9a0c803
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat1_y_net,
      d1 => register2_q_net_x6,
      y => logical1_y_net
    );

  map_rom: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 12,
      c_address_width_b => 12,
      c_width_a => 9,
      c_width_b => 9,
      core_name0 => "bmg_72_30fab105208816ae",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x57,
      a_clk => clk_1_sg_x57,
      addra => concat2_y_net,
      addrb => concat3_y_net,
      b_ce => ce_1_sg_x57,
      b_clk => clk_1_sg_x57,
      dina => constant8_op_net,
      dinb => constant8_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant9_op_net,
      web(0) => constant9_op_net,
      douta => map_rom_douta_net_x1,
      doutb => map_rom_doutb_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Puncturing/Rate 1/2"

entity x2_entity_63e54e2fbc is
  port (
    ind_inc: out std_logic_vector(1 downto 0); 
    skip_a: out std_logic
  );
end x2_entity_63e54e2fbc;

architecture structural of x2_entity_63e54e2fbc is
  signal constant2_op_net_x0: std_logic;
  signal constant3_op_net_x0: std_logic_vector(1 downto 0);

begin
  ind_inc <= constant3_op_net_x0;
  skip_a <= constant2_op_net_x0;

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net_x0
    );

  constant3: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Puncturing/Rate 2/3"

entity x3_entity_e9b5af3b14 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    ind_inc: out std_logic_vector(1 downto 0); 
    skip_a: out std_logic; 
    skip_b: out std_logic
  );
end x3_entity_e9b5af3b14;

architecture structural of x3_entity_e9b5af3b14 is
  signal ce_1_sg_x58: std_logic;
  signal clk_1_sg_x58: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net_x0: std_logic;
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal delay3_q_net_x2: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal mux3_y_net_x0: std_logic_vector(1 downto 0);
  signal relational_op_net_x0: std_logic;
  signal x0_1_op_net: std_logic;

begin
  ce_1_sg_x58 <= ce_1;
  clk_1_sg_x58 <= clk_1;
  delay3_q_net_x2 <= en;
  logical2_y_net_x1 <= rst;
  ind_inc <= mux3_y_net_x0;
  skip_a <= constant2_op_net_x0;
  skip_b <= relational_op_net_x0;

  constant1: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net_x0
    );

  constant3: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  mux3: entity work.mux_2a63ac73aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant3_op_net,
      d1 => constant4_op_net,
      sel(0) => relational_op_net_x0,
      y => mux3_y_net_x0
    );

  relational: entity work.relational_194eb61c1b
    port map (
      a(0) => x0_1_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net_x0
    );

  x0_1: entity work.counter_caa2b01eef
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      en(0) => delay3_q_net_x2,
      rst(0) => logical2_y_net_x1,
      op(0) => x0_1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Puncturing/Rate 3/4"

entity x4_entity_e63825ace3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    ind_inc: out std_logic_vector(1 downto 0); 
    skip_a: out std_logic; 
    skip_b: out std_logic
  );
end x4_entity_e63825ace3;

architecture structural of x4_entity_e63825ace3 is
  signal ce_1_sg_x59: std_logic;
  signal clk_1_sg_x59: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal constant7_op_net: std_logic_vector(1 downto 0);
  signal delay3_q_net_x3: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal mux3_y_net_x0: std_logic_vector(1 downto 0);
  signal relational2_op_net_x0: std_logic;
  signal relational_op_net_x0: std_logic;
  signal x0_2_op_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x59 <= ce_1;
  clk_1_sg_x59 <= clk_1;
  delay3_q_net_x3 <= en;
  logical2_y_net_x2 <= rst;
  ind_inc <= mux3_y_net_x0;
  skip_a <= relational_op_net_x0;
  skip_b <= relational2_op_net_x0;

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => relational2_op_net_x0,
      in1(0) => relational_op_net_x0,
      y => concat_y_net
    );

  constant1: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant7: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net
    );

  mux3: entity work.mux_78aa6a36ae
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant3_op_net,
      d1 => constant4_op_net,
      d2 => constant7_op_net,
      sel => concat_y_net,
      y => mux3_y_net_x0
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => x0_2_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net_x0
    );

  relational2: entity work.relational_f52e6abf76
    port map (
      a => x0_2_op_net,
      b(0) => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net_x0
    );

  x0_2: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 2,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_6454489cfe866515",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      en(0) => delay3_q_net_x3,
      rst(0) => logical2_y_net_x2,
      op => x0_2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Puncturing/Rate 5/6"

entity x6_entity_01983fe4c9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    ind_inc: out std_logic_vector(1 downto 0); 
    skip_a: out std_logic; 
    skip_b: out std_logic
  );
end x6_entity_01983fe4c9;

architecture structural of x6_entity_01983fe4c9 is
  signal ce_1_sg_x60: std_logic;
  signal clk_1_sg_x60: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal constant5_op_net: std_logic_vector(1 downto 0);
  signal constant6_op_net: std_logic_vector(2 downto 0);
  signal constant7_op_net: std_logic_vector(1 downto 0);
  signal delay3_q_net_x4: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net_x3: std_logic;
  signal logical_y_net_x0: std_logic;
  signal mux3_y_net_x0: std_logic_vector(1 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational_op_net: std_logic;
  signal x0_4_op_net: std_logic_vector(2 downto 0);

begin
  ce_1_sg_x60 <= ce_1;
  clk_1_sg_x60 <= clk_1;
  delay3_q_net_x4 <= en;
  logical2_y_net_x3 <= rst;
  ind_inc <= mux3_y_net_x0;
  skip_a <= logical_y_net_x0;
  skip_b <= logical1_y_net_x0;

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => logical1_y_net_x0,
      in1(0) => logical_y_net_x0,
      y => concat_y_net
    );

  constant1: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  constant7: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational_op_net,
      d1(0) => relational2_op_net,
      y(0) => logical_y_net_x0
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net,
      d1(0) => relational3_op_net,
      y(0) => logical1_y_net_x0
    );

  mux3: entity work.mux_78aa6a36ae
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant3_op_net,
      d1 => constant4_op_net,
      d2 => constant7_op_net,
      sel => concat_y_net,
      y => mux3_y_net_x0
    );

  relational: entity work.relational_706b9eb7ce
    port map (
      a => x0_4_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_706b9eb7ce
    port map (
      a => x0_4_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_8fc7f5539b
    port map (
      a => x0_4_op_net,
      b => constant6_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_706b9eb7ce
    port map (
      a => x0_4_op_net,
      b => constant5_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  x0_4: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 4,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_bcc28bfecf25caff",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 3
    )
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      en(0) => delay3_q_net_x4,
      rst(0) => logical2_y_net_x3,
      op => x0_4_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/Puncturing"

entity puncturing_entity_bd1c34b968 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    code_rate: in std_logic_vector(1 downto 0); 
    en: in std_logic; 
    reset: in std_logic; 
    index_inc: out std_logic_vector(1 downto 0); 
    wr_a: out std_logic; 
    wr_b: out std_logic
  );
end puncturing_entity_bd1c34b968;

architecture structural of puncturing_entity_bd1c34b968 is
  signal ce_1_sg_x61: std_logic;
  signal clk_1_sg_x61: std_logic;
  signal constant2_op_net_x0: std_logic;
  signal constant2_op_net_x1: std_logic;
  signal constant3_op_net_x0: std_logic_vector(1 downto 0);
  signal delay3_q_net_x5: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x4: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x1: std_logic;
  signal mux1_y_net: std_logic;
  signal mux2_y_net_x0: std_logic_vector(1 downto 0);
  signal mux3_y_net: std_logic;
  signal mux3_y_net_x0: std_logic_vector(1 downto 0);
  signal mux3_y_net_x1: std_logic_vector(1 downto 0);
  signal mux3_y_net_x2: std_logic_vector(1 downto 0);
  signal mux4_y_net_x1: std_logic_vector(1 downto 0);
  signal relational2_op_net_x0: std_logic;
  signal relational_op_net_x0: std_logic;
  signal relational_op_net_x1: std_logic;

begin
  ce_1_sg_x61 <= ce_1;
  clk_1_sg_x61 <= clk_1;
  mux2_y_net_x0 <= code_rate;
  delay3_q_net_x5 <= en;
  logical2_y_net_x4 <= reset;
  index_inc <= mux4_y_net_x1;
  wr_a <= logical_y_net_x1;
  wr_b <= logical1_y_net_x1;

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      ip(0) => mux3_y_net,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      ip(0) => mux1_y_net,
      op(0) => inverter1_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => delay3_q_net_x5,
      y(0) => logical_y_net_x1
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter1_op_net,
      d1(0) => delay3_q_net_x5,
      y(0) => logical1_y_net_x1
    );

  mux1: entity work.mux_cdffdf53c9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => constant2_op_net_x0,
      d1(0) => relational_op_net_x0,
      d2(0) => relational2_op_net_x0,
      d3(0) => logical1_y_net_x0,
      sel => mux2_y_net_x0,
      y(0) => mux1_y_net
    );

  mux3: entity work.mux_cdffdf53c9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => constant2_op_net_x0,
      d1(0) => constant2_op_net_x1,
      d2(0) => relational_op_net_x1,
      d3(0) => logical_y_net_x0,
      sel => mux2_y_net_x0,
      y(0) => mux3_y_net
    );

  mux4: entity work.mux_1a0db76efe
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant3_op_net_x0,
      d1 => mux3_y_net_x0,
      d2 => mux3_y_net_x1,
      d3 => mux3_y_net_x2,
      sel => mux2_y_net_x0,
      y => mux4_y_net_x1
    );

  x2_63e54e2fbc: entity work.x2_entity_63e54e2fbc
    port map (
      ind_inc => constant3_op_net_x0,
      skip_a => constant2_op_net_x0
    );

  x3_e9b5af3b14: entity work.x3_entity_e9b5af3b14
    port map (
      ce_1 => ce_1_sg_x61,
      clk_1 => clk_1_sg_x61,
      en => delay3_q_net_x5,
      rst => logical2_y_net_x4,
      ind_inc => mux3_y_net_x0,
      skip_a => constant2_op_net_x1,
      skip_b => relational_op_net_x0
    );

  x4_e63825ace3: entity work.x4_entity_e63825ace3
    port map (
      ce_1 => ce_1_sg_x61,
      clk_1 => clk_1_sg_x61,
      en => delay3_q_net_x5,
      rst => logical2_y_net_x4,
      ind_inc => mux3_y_net_x1,
      skip_a => relational_op_net_x1,
      skip_b => relational2_op_net_x0
    );

  x6_01983fe4c9: entity work.x6_entity_01983fe4c9
    port map (
      ce_1 => ce_1_sg_x61,
      clk_1 => clk_1_sg_x61,
      en => delay3_q_net_x5,
      rst => logical2_y_net_x4,
      ind_inc => mux3_y_net_x2,
      skip_a => logical_y_net_x0,
      skip_b => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing/negedge"

entity negedge_entity_02af90a306 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end negedge_entity_02af90a306;

architecture structural of negedge_entity_02af90a306 is
  signal ce_1_sg_x62: std_logic;
  signal clk_1_sg_x62: std_logic;
  signal delay3_q_net_x6: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;

begin
  ce_1_sg_x62 <= ce_1;
  clk_1_sg_x62 <= clk_1;
  delay3_q_net_x6 <= d;
  q <= logical1_y_net_x0;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x62,
      clk => clk_1_sg_x62,
      d(0) => delay3_q_net_x6,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x62,
      clk => clk_1_sg_x62,
      clr => '0',
      ip(0) => delay3_q_net_x6,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Interleaver Ctrl & Puncturing"

entity \interleaver_ctrl___puncturing_entity_e6d742099d\ is
  port (
    base_rate: in std_logic; 
    bits_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ofdm_tx_data_code_rate: in std_logic_vector(1 downto 0); 
    pkt_data: in std_logic_vector(1 downto 0); 
    slice1: in std_logic; 
    tx_reset: in std_logic; 
    addr_a: out std_logic_vector(8 downto 0); 
    addr_b: out std_logic_vector(8 downto 0); 
    wr_a: out std_logic; 
    wr_b: out std_logic
  );
end \interleaver_ctrl___puncturing_entity_e6d742099d\;

architecture structural of \interleaver_ctrl___puncturing_entity_e6d742099d\ is
  signal accumulator_q_net_x1: std_logic_vector(8 downto 0);
  signal addsub_s_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x63: std_logic;
  signal clk_1_sg_x63: std_logic;
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x3: std_logic;
  signal delay2_q_net_x3: std_logic;
  signal delay3_q_net_x7: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x4: std_logic;
  signal logical_y_net_x1: std_logic;
  signal logical_y_net_x30: std_logic;
  signal map_rom_douta_net_x2: std_logic_vector(8 downto 0);
  signal map_rom_doutb_net_x2: std_logic_vector(8 downto 0);
  signal mcode_load_base_rate_net_x1: std_logic;
  signal mux2_y_net_x0: std_logic_vector(1 downto 0);
  signal mux4_y_net_x1: std_logic_vector(1 downto 0);
  signal register2_q_net_x7: std_logic_vector(1 downto 0);
  signal register3_q_net_x2: std_logic_vector(1 downto 0);
  signal slice1_y_net_x10: std_logic;

begin
  mcode_load_base_rate_net_x1 <= base_rate;
  delay3_q_net_x7 <= bits_tvalid;
  ce_1_sg_x63 <= ce_1;
  clk_1_sg_x63 <= clk_1;
  register3_q_net_x2 <= ofdm_tx_data_code_rate;
  register2_q_net_x7 <= pkt_data;
  slice1_y_net_x10 <= slice1;
  logical_y_net_x30 <= tx_reset;
  addr_a <= map_rom_douta_net_x2;
  addr_b <= map_rom_doutb_net_x2;
  wr_a <= delay1_q_net_x3;
  wr_b <= delay2_q_net_x3;

  bit_index_calc_ec83e953ec: entity work.bit_index_calc_entity_ec83e953ec
    port map (
      ce_1 => ce_1_sg_x63,
      clk_1 => clk_1_sg_x63,
      en => delay3_q_net_x7,
      inc => mux4_y_net_x1,
      rst => logical2_y_net_x4,
      ind_a => accumulator_q_net_x1,
      ind_b => addsub_s_net_x1
    );

  constant2: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d(0) => logical_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x3
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d(0) => logical1_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x3
    );

  interleave_mapping_48a573e6d3: entity work.interleave_mapping_entity_48a573e6d3
    port map (
      base_rate_sym => mcode_load_base_rate_net_x1,
      ce_1 => ce_1_sg_x63,
      clk_1 => clk_1_sg_x63,
      ind_a => accumulator_q_net_x1,
      ind_b => addsub_s_net_x1,
      ofdm_tx_data_mod_sel => register2_q_net_x7,
      tx_phy_mode_11n => slice1_y_net_x10,
      addr_a => map_rom_douta_net_x2,
      addr_b => map_rom_doutb_net_x2
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x30,
      d1(0) => logical1_y_net_x0,
      y(0) => logical2_y_net_x4
    );

  mux2: entity work.mux_2a63ac73aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register3_q_net_x2,
      d1 => constant2_op_net,
      sel(0) => mcode_load_base_rate_net_x1,
      y => mux2_y_net_x0
    );

  negedge_02af90a306: entity work.negedge_entity_02af90a306
    port map (
      ce_1 => ce_1_sg_x63,
      clk_1 => clk_1_sg_x63,
      d => delay3_q_net_x7,
      q => logical1_y_net_x0
    );

  puncturing_bd1c34b968: entity work.puncturing_entity_bd1c34b968
    port map (
      ce_1 => ce_1_sg_x63,
      clk_1 => clk_1_sg_x63,
      code_rate => mux2_y_net_x0,
      en => delay3_q_net_x7,
      reset => logical2_y_net_x4,
      index_inc => mux4_y_net_x1,
      wr_a => logical_y_net_x1,
      wr_b => logical1_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave/Mem Sel"

entity mem_sel_entity_0052fdd6ac is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    tx_reset: in std_logic; 
    rd: out std_logic; 
    wr: out std_logic
  );
end mem_sel_entity_0052fdd6ac;

architecture structural of mem_sel_entity_0052fdd6ac is
  signal ce_1_sg_x65: std_logic;
  signal clk_1_sg_x65: std_logic;
  signal delay4_q_net_x0: std_logic;
  signal inverter_op_net_x1: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x31: std_logic;
  signal register2_q_net_x2: std_logic;

begin
  ce_1_sg_x65 <= ce_1;
  clk_1_sg_x65 <= clk_1;
  delay4_q_net_x0 <= en;
  logical_y_net_x31 <= tx_reset;
  rd <= register2_q_net_x2;
  wr <= inverter_op_net_x1;

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x65,
      clk => clk_1_sg_x65,
      clr => '0',
      ip(0) => register2_q_net_x2,
      op(0) => inverter_op_net_x1
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net_x1,
      d1(0) => delay4_q_net_x0,
      y(0) => logical_y_net_x0
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay4_q_net_x0,
      d1(0) => register2_q_net_x2,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net,
      d1(0) => logical_y_net_x31,
      y(0) => logical2_y_net_x0
    );

  s_r_latch1_1b9e9bb936: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x65,
      clk_1 => clk_1_sg_x65,
      r => logical2_y_net_x0,
      s => logical_y_net_x0,
      q => register2_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen/Puncture & Interleave"

entity \puncture___interleave_entity_fa36f44c5c\ is
  port (
    bit_a: in std_logic; 
    bit_b: in std_logic; 
    bits_tlast: in std_logic; 
    bits_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_sym_ind: in std_logic_vector(5 downto 0); 
    logical: in std_logic; 
    pkt_data: in std_logic_vector(1 downto 0); 
    pkt_data_x0: in std_logic_vector(1 downto 0); 
    slice1: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    sc_bits: out std_logic_vector(7 downto 0); 
    sym_bits_rdy: out std_logic; 
    sym_cfg_x0: out std_logic_vector(17 downto 0)
  );
end \puncture___interleave_entity_fa36f44c5c\;

architecture structural of \puncture___interleave_entity_fa36f44c5c\ is
  signal a_xor_y_net_x1: std_logic;
  signal b_xor_y_net_x1: std_logic;
  signal ce_1_sg_x66: std_logic;
  signal clk_1_sg_x66: std_logic;
  signal delay1_q_net_x1: std_logic;
  signal delay1_q_net_x3: std_logic;
  signal delay1_q_net_x4: std_logic_vector(17 downto 0);
  signal delay2_q_net_x1: std_logic;
  signal delay2_q_net_x3: std_logic;
  signal delay2_q_net_x4: std_logic;
  signal delay3_q_net: std_logic_vector(17 downto 0);
  signal delay3_q_net_x8: std_logic;
  signal delay4_q_net_x0: std_logic;
  signal delay5_q_net_x4: std_logic;
  signal delay6_q_net_x2: std_logic_vector(17 downto 0);
  signal inverter_op_net_x1: std_logic;
  signal logical_y_net_x32: std_logic;
  signal map_rom_douta_net_x2: std_logic_vector(8 downto 0);
  signal map_rom_doutb_net_x2: std_logic_vector(8 downto 0);
  signal mcode_load_base_rate_net_x1: std_logic;
  signal mux1_y_net_x7: std_logic_vector(7 downto 0);
  signal register2_q_net_x2: std_logic;
  signal register2_q_net_x8: std_logic_vector(1 downto 0);
  signal register3_q_net_x3: std_logic_vector(1 downto 0);
  signal slice1_y_net_x11: std_logic;
  signal slice_y_net_x4: std_logic_vector(5 downto 0);

begin
  a_xor_y_net_x1 <= bit_a;
  b_xor_y_net_x1 <= bit_b;
  delay2_q_net_x4 <= bits_tlast;
  delay3_q_net_x8 <= bits_tvalid;
  ce_1_sg_x66 <= ce_1;
  clk_1_sg_x66 <= clk_1;
  slice_y_net_x4 <= data_sym_ind;
  logical_y_net_x32 <= logical;
  register2_q_net_x8 <= pkt_data;
  register3_q_net_x3 <= pkt_data_x0;
  slice1_y_net_x11 <= slice1;
  delay1_q_net_x4 <= sym_cfg;
  sc_bits <= mux1_y_net_x7;
  sym_bits_rdy <= delay5_q_net_x4;
  sym_cfg_x0 <= delay6_q_net_x2;

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d(0) => a_xor_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x1
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d(0) => b_xor_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x1
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d => delay1_q_net_x4,
      en => '1',
      rst => '1',
      q => delay3_q_net
    );

  delay4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d(0) => delay2_q_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay4_q_net_x0
    );

  delay5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d(0) => delay4_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay5_q_net_x4
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 18
    )
    port map (
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      d => delay3_q_net,
      en => delay2_q_net_x3,
      rst => '1',
      q => delay6_q_net_x2
    );

  interleave_ram_42ac73a366: entity work.interleave_ram_entity_42ac73a366
    port map (
      bit_a => delay1_q_net_x1,
      bit_addr_a => map_rom_douta_net_x2,
      bit_addr_b => map_rom_doutb_net_x2,
      bit_b => delay2_q_net_x1,
      ce_1 => ce_1_sg_x66,
      clk_1 => clk_1_sg_x66,
      rd_addr => slice_y_net_x4,
      rd_mem_sel => register2_q_net_x2,
      wr_a => delay1_q_net_x3,
      wr_b => delay2_q_net_x3,
      wr_mem_sel => inverter_op_net_x1,
      sc_bits => mux1_y_net_x7
    );

  interleaver_ctrl_puncturing_e6d742099d: entity work.\interleaver_ctrl___puncturing_entity_e6d742099d\
    port map (
      base_rate => mcode_load_base_rate_net_x1,
      bits_tvalid => delay3_q_net_x8,
      ce_1 => ce_1_sg_x66,
      clk_1 => clk_1_sg_x66,
      ofdm_tx_data_code_rate => register3_q_net_x3,
      pkt_data => register2_q_net_x8,
      slice1 => slice1_y_net_x11,
      tx_reset => logical_y_net_x32,
      addr_a => map_rom_douta_net_x2,
      addr_b => map_rom_doutb_net_x2,
      wr_a => delay1_q_net_x3,
      wr_b => delay2_q_net_x3
    );

  mcode: entity work.mcode_block_00412594a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      sym_cfg => delay1_q_net_x4,
      load_base_rate(0) => mcode_load_base_rate_net_x1
    );

  mem_sel_0052fdd6ac: entity work.mem_sel_entity_0052fdd6ac
    port map (
      ce_1 => ce_1_sg_x66,
      clk_1 => clk_1_sg_x66,
      en => delay4_q_net_x0,
      tx_reset => logical_y_net_x32,
      rd => register2_q_net_x2,
      wr => inverter_op_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/PSDU Syms Gen"

entity psdu_syms_gen_entity_1449f55c9b is
  port (
    bram_din: in std_logic_vector(63 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    iq_fifo_tready: in std_logic; 
    logical: in std_logic; 
    logical3: in std_logic; 
    mux: in std_logic_vector(3 downto 0); 
    register16: in std_logic_vector(7 downto 0); 
    register2: in std_logic; 
    register8: in std_logic_vector(7 downto 0); 
    slice: in std_logic; 
    slice1: in std_logic; 
    start_sym: in std_logic; 
    sym_cfg: in std_logic_vector(17 downto 0); 
    data_done: out std_logic; 
    iq_stream: out std_logic_vector(11 downto 0); 
    modulate: out std_logic; 
    modulate_x0: out std_logic; 
    modulate_x1: out std_logic_vector(11 downto 0); 
    pkt_data: out std_logic_vector(31 downto 0); 
    pkt_data_x0: out std_logic; 
    pkt_data_x1: out std_logic; 
    pkt_data_x2: out std_logic_vector(63 downto 0); 
    pkt_data_x3: out std_logic_vector(7 downto 0); 
    pkt_data_x4: out std_logic; 
    sym_cfg_x0: out std_logic_vector(17 downto 0)
  );
end psdu_syms_gen_entity_1449f55c9b;

architecture structural of psdu_syms_gen_entity_1449f55c9b is
  signal a_xor_y_net_x1: std_logic;
  signal axi_fifo_s_axis_tready_net_x5: std_logic;
  signal b_xor_y_net_x1: std_logic;
  signal bit_in_byte_y_net_x3: std_logic_vector(2 downto 0);
  signal bram_din_net_x3: std_logic_vector(63 downto 0);
  signal bytes_y_net_x4: std_logic_vector(11 downto 0);
  signal ce_1_sg_x67: std_logic;
  signal clk_1_sg_x67: std_logic;
  signal concat_y_net_x3: std_logic_vector(31 downto 0);
  signal concat_y_net_x7: std_logic_vector(17 downto 0);
  signal constant1_op_net_x3: std_logic;
  signal constant2_op_net_x3: std_logic;
  signal constant7_op_net_x3: std_logic_vector(63 downto 0);
  signal constant8_op_net_x3: std_logic_vector(7 downto 0);
  signal delay1_q_net_x3: std_logic;
  signal delay1_q_net_x4: std_logic_vector(17 downto 0);
  signal delay2_q_net_x3: std_logic;
  signal delay2_q_net_x4: std_logic;
  signal delay3_q_net_x8: std_logic;
  signal delay5_q_net_x4: std_logic;
  signal delay6_q_net_x2: std_logic_vector(17 downto 0);
  signal delay8_q_net_x1: std_logic_vector(17 downto 0);
  signal delay9_q_net_x3: std_logic;
  signal delay_q_net_x8: std_logic;
  signal delay_q_net_x9: std_logic_vector(17 downto 0);
  signal logical1_y_net_x2: std_logic;
  signal logical3_y_net_x6: std_logic;
  signal logical4_y_net_x4: std_logic;
  signal logical4_y_net_x7: std_logic;
  signal logical4_y_net_x8: std_logic;
  signal logical5_y_net_x2: std_logic;
  signal logical_y_net_x2: std_logic;
  signal logical_y_net_x33: std_logic;
  signal mux1_y_net_x7: std_logic_vector(7 downto 0);
  signal mux3_y_net_x2: std_logic_vector(11 downto 0);
  signal mux4_y_net_x2: std_logic_vector(11 downto 0);
  signal mux_y_net_x12: std_logic_vector(3 downto 0);
  signal register16_q_net_x2: std_logic_vector(7 downto 0);
  signal register1_q_net_x3: std_logic_vector(9 downto 0);
  signal register2_q_net_x5: std_logic;
  signal register2_q_net_x8: std_logic_vector(1 downto 0);
  signal register3_q_net_x3: std_logic_vector(1 downto 0);
  signal register8_q_net_x8: std_logic_vector(7 downto 0);
  signal slice1_y_net_x12: std_logic;
  signal slice_y_net_x4: std_logic_vector(5 downto 0);
  signal slice_y_net_x5: std_logic;

begin
  bram_din_net_x3 <= bram_din;
  ce_1_sg_x67 <= ce_1;
  clk_1_sg_x67 <= clk_1;
  axi_fifo_s_axis_tready_net_x5 <= iq_fifo_tready;
  logical_y_net_x33 <= logical;
  logical3_y_net_x6 <= logical3;
  mux_y_net_x12 <= mux;
  register16_q_net_x2 <= register16;
  register2_q_net_x5 <= register2;
  register8_q_net_x8 <= register8;
  slice_y_net_x5 <= slice;
  slice1_y_net_x12 <= slice1;
  logical4_y_net_x7 <= start_sym;
  concat_y_net_x7 <= sym_cfg;
  data_done <= delay9_q_net_x3;
  iq_stream <= mux3_y_net_x2;
  modulate <= delay_q_net_x8;
  modulate_x0 <= delay1_q_net_x3;
  modulate_x1 <= mux4_y_net_x2;
  pkt_data <= concat_y_net_x3;
  pkt_data_x0 <= constant1_op_net_x3;
  pkt_data_x1 <= constant2_op_net_x3;
  pkt_data_x2 <= constant7_op_net_x3;
  pkt_data_x3 <= constant8_op_net_x3;
  pkt_data_x4 <= logical4_y_net_x8;
  sym_cfg_x0 <= delay_q_net_x9;

  convolutional_encoder_c777b8e511: entity work.convolutional_encoder_entity_c777b8e511
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      sym_cfg => delay8_q_net_x1,
      tx_bit => logical_y_net_x2,
      tx_bit_tlast => logical1_y_net_x2,
      tx_bit_tvalid => delay2_q_net_x3,
      tx_reset => logical_y_net_x33,
      enc_bit_a => a_xor_y_net_x1,
      enc_bit_b => b_xor_y_net_x1,
      enc_bits_tlast => delay2_q_net_x4,
      enc_bits_tvalid => delay3_q_net_x8,
      sym_cfg_x0 => delay1_q_net_x4
    );

  index_gen_b965cbdf90: entity work.index_gen_entity_b965cbdf90
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      logical => logical_y_net_x33,
      register1 => register1_q_net_x3,
      start_sym => logical4_y_net_x7,
      sym_cfg => concat_y_net_x7,
      bit_sel => bit_in_byte_y_net_x3,
      bit_sel_valid => logical4_y_net_x4,
      byte_ind => bytes_y_net_x4,
      byte_ind_valid => logical5_y_net_x2
    );

  modulate_324fd14050: entity work.modulate_entity_324fd14050
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      iq_fifo_tready => axi_fifo_s_axis_tready_net_x5,
      logical => logical_y_net_x33,
      ofdm_tx_data_mod_sel => register2_q_net_x8,
      register8 => register8_q_net_x8,
      sc_bits => mux1_y_net_x7,
      slice1 => slice1_y_net_x12,
      sym_bits_rdy => delay5_q_net_x4,
      sym_cfg => delay6_q_net_x2,
      data_sym_ind => slice_y_net_x4,
      i => mux3_y_net_x2,
      iq_tlast => delay1_q_net_x3,
      iq_tvalid => delay_q_net_x8,
      q => mux4_y_net_x2,
      sym_cfg_x0 => delay_q_net_x9
    );

  pkt_data_6db78f9ff0: entity work.pkt_data_entity_6db78f9ff0
    port map (
      bit_sel => bit_in_byte_y_net_x3,
      bit_sel_valid => logical4_y_net_x4,
      bram_din => bram_din_net_x3,
      byte_ind => bytes_y_net_x4,
      byte_ind_valid => logical5_y_net_x2,
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      logical => logical_y_net_x33,
      logical3 => logical3_y_net_x6,
      mux => mux_y_net_x12,
      register16 => register16_q_net_x2,
      register2 => register2_q_net_x5,
      slice => slice_y_net_x5,
      slice1 => slice1_y_net_x12,
      sym_cfg => concat_y_net_x7,
      bram_if_64b => concat_y_net_x3,
      bram_if_64b_x0 => constant1_op_net_x3,
      bram_if_64b_x1 => constant2_op_net_x3,
      bram_if_64b_x2 => constant7_op_net_x3,
      bram_if_64b_x3 => constant8_op_net_x3,
      data_done => delay9_q_net_x3,
      signal_ht_sig_decode => register1_q_net_x3,
      signal_ht_sig_decode_x0 => register2_q_net_x8,
      signal_ht_sig_decode_x1 => register3_q_net_x3,
      sym_cfg_x0 => delay8_q_net_x1,
      tx_bit => logical_y_net_x2,
      tx_bit_tlast => logical1_y_net_x2,
      tx_bit_tvalid => delay2_q_net_x3,
      tx_sig_decode_error => logical4_y_net_x8
    );

  puncture_interleave_fa36f44c5c: entity work.\puncture___interleave_entity_fa36f44c5c\
    port map (
      bit_a => a_xor_y_net_x1,
      bit_b => b_xor_y_net_x1,
      bits_tlast => delay2_q_net_x4,
      bits_tvalid => delay3_q_net_x8,
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      data_sym_ind => slice_y_net_x4,
      logical => logical_y_net_x33,
      pkt_data => register2_q_net_x8,
      pkt_data_x0 => register3_q_net_x3,
      slice1 => slice1_y_net_x12,
      sym_cfg => delay1_q_net_x4,
      sc_bits => mux1_y_net_x7,
      sym_bits_rdy => delay5_q_net_x4,
      sym_cfg_x0 => delay6_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/DAC Outputs/Ant Enables"

entity ant_enables_entity_b219a59ac1 is
  port (
    mac_tx_ant_mask: in std_logic_vector(3 downto 0); 
    regtx_anta_tx_en: in std_logic; 
    regtx_antb_tx_en: in std_logic; 
    regtx_antc_tx_en: in std_logic; 
    regtx_antd_tx_en: in std_logic; 
    regtx_use_mac_ant_masks: in std_logic; 
    a_en: out std_logic; 
    b_en: out std_logic; 
    c_en: out std_logic; 
    d_en: out std_logic
  );
end ant_enables_entity_b219a59ac1;

architecture structural of ant_enables_entity_b219a59ac1 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net_x0: std_logic;
  signal logical5_y_net: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical7_y_net: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal register1_q_net_x0: std_logic_vector(3 downto 0);
  signal register23_q_net_x0: std_logic;
  signal register3_q_net_x0: std_logic;
  signal register4_q_net_x0: std_logic;
  signal register5_q_net_x0: std_logic;
  signal register6_q_net_x0: std_logic;

begin
  register1_q_net_x0 <= mac_tx_ant_mask;
  register3_q_net_x0 <= regtx_anta_tx_en;
  register4_q_net_x0 <= regtx_antb_tx_en;
  register5_q_net_x0 <= regtx_antc_tx_en;
  register6_q_net_x0 <= regtx_antd_tx_en;
  register23_q_net_x0 <= regtx_use_mac_ant_masks;
  a_en <= logical2_y_net_x0;
  b_en <= logical4_y_net_x0;
  c_en <= logical6_y_net_x0;
  d_en <= logical8_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x0,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x0,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x0,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x0,
      y(0) => b3_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b0_y_net,
      d1(0) => register23_q_net_x0,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register3_q_net_x0,
      d1(0) => logical1_y_net,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b1_y_net,
      d1(0) => register23_q_net_x0,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register4_q_net_x0,
      d1(0) => logical3_y_net,
      y(0) => logical4_y_net_x0
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b2_y_net,
      d1(0) => register23_q_net_x0,
      y(0) => logical5_y_net
    );

  logical6: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register5_q_net_x0,
      d1(0) => logical5_y_net,
      y(0) => logical6_y_net_x0
    );

  logical7: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b3_y_net,
      d1(0) => register23_q_net_x0,
      y(0) => logical7_y_net
    );

  logical8: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register6_q_net_x0,
      d1(0) => logical7_y_net,
      y(0) => logical8_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/DAC Outputs"

entity dac_outputs_entity_fec48642b9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    i: in std_logic_vector(11 downto 0); 
    q: in std_logic_vector(11 downto 0); 
    register1_x0: in std_logic_vector(3 downto 0); 
    register23: in std_logic; 
    register3_x0: in std_logic; 
    register4_x0: in std_logic; 
    register5_x0: in std_logic; 
    register6_x0: in std_logic; 
    register1_x1: out std_logic_vector(11 downto 0); 
    register2_x0: out std_logic_vector(11 downto 0); 
    register3_x1: out std_logic_vector(11 downto 0); 
    register4_x1: out std_logic_vector(11 downto 0); 
    register5_x1: out std_logic_vector(11 downto 0); 
    register6_x1: out std_logic_vector(11 downto 0); 
    register7_x0: out std_logic_vector(11 downto 0); 
    register_x1: out std_logic_vector(11 downto 0)
  );
end dac_outputs_entity_fec48642b9;

architecture structural of dac_outputs_entity_fec48642b9 is
  signal ce_1_sg_x68: std_logic;
  signal clk_1_sg_x68: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal inverter4_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net_x0: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mult1_p_net_x0: std_logic_vector(11 downto 0);
  signal mult_p_net_x0: std_logic_vector(11 downto 0);
  signal register10_q_net: std_logic_vector(11 downto 0);
  signal register1_q_net_x1: std_logic_vector(3 downto 0);
  signal register1_q_net_x2: std_logic_vector(11 downto 0);
  signal register23_q_net_x1: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x2: std_logic_vector(11 downto 0);
  signal register3_q_net_x1: std_logic;
  signal register3_q_net_x2: std_logic_vector(11 downto 0);
  signal register4_q_net_x1: std_logic;
  signal register4_q_net_x2: std_logic_vector(11 downto 0);
  signal register5_q_net_x1: std_logic;
  signal register5_q_net_x2: std_logic_vector(11 downto 0);
  signal register6_q_net_x1: std_logic;
  signal register6_q_net_x2: std_logic_vector(11 downto 0);
  signal register7_q_net_x0: std_logic_vector(11 downto 0);
  signal register8_q_net: std_logic_vector(11 downto 0);
  signal register9_q_net: std_logic;
  signal register_q_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x68 <= ce_1;
  clk_1_sg_x68 <= clk_1;
  register2_q_net_x1 <= en;
  mult_p_net_x0 <= i;
  mult1_p_net_x0 <= q;
  register1_q_net_x1 <= register1_x0;
  register23_q_net_x1 <= register23;
  register3_q_net_x1 <= register3_x0;
  register4_q_net_x1 <= register4_x0;
  register5_q_net_x1 <= register5_x0;
  register6_q_net_x1 <= register6_x0;
  register1_x1 <= register1_q_net_x2;
  register2_x0 <= register2_q_net_x2;
  register3_x1 <= register3_q_net_x2;
  register4_x1 <= register4_q_net_x2;
  register5_x1 <= register5_q_net_x2;
  register6_x1 <= register6_q_net_x2;
  register7_x0 <= register7_q_net_x0;
  register_x1 <= register_q_net_x0;

  ant_enables_b219a59ac1: entity work.ant_enables_entity_b219a59ac1
    port map (
      mac_tx_ant_mask => register1_q_net_x1,
      regtx_anta_tx_en => register3_q_net_x1,
      regtx_antb_tx_en => register4_q_net_x1,
      regtx_antc_tx_en => register5_q_net_x1,
      regtx_antd_tx_en => register6_q_net_x1,
      regtx_use_mac_ant_masks => register23_q_net_x1,
      a_en => logical2_y_net_x0,
      b_en => logical4_y_net_x0,
      c_en => logical6_y_net_x0,
      d_en => logical8_y_net_x0
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      clr => '0',
      ip(0) => logical_y_net,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      clr => '0',
      ip(0) => logical1_y_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      clr => '0',
      ip(0) => logical2_y_net,
      op(0) => inverter3_op_net
    );

  inverter4: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      clr => '0',
      ip(0) => logical3_y_net,
      op(0) => inverter4_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register9_q_net,
      d1(0) => logical2_y_net_x0,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register9_q_net,
      d1(0) => logical4_y_net_x0,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register9_q_net,
      d1(0) => logical6_y_net_x0,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register9_q_net,
      d1(0) => logical8_y_net_x0,
      y(0) => logical3_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register10_q_net,
      en => "1",
      rst(0) => inverter1_op_net,
      q => register1_q_net_x2
    );

  register10: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => mult1_p_net_x0,
      en => "1",
      rst => "0",
      q => register10_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register8_q_net,
      en => "1",
      rst(0) => inverter2_op_net,
      q => register2_q_net_x2
    );

  register3: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register10_q_net,
      en => "1",
      rst(0) => inverter2_op_net,
      q => register3_q_net_x2
    );

  register4: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register8_q_net,
      en => "1",
      rst(0) => inverter3_op_net,
      q => register4_q_net_x2
    );

  register5: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register10_q_net,
      en => "1",
      rst(0) => inverter3_op_net,
      q => register5_q_net_x2
    );

  register6: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register8_q_net,
      en => "1",
      rst(0) => inverter4_op_net,
      q => register6_q_net_x2
    );

  register7: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register10_q_net,
      en => "1",
      rst(0) => inverter4_op_net,
      q => register7_q_net_x0
    );

  register8: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => mult_p_net_x0,
      en => "1",
      rst => "0",
      q => register8_q_net
    );

  register9: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d(0) => register2_q_net_x1,
      en => "1",
      rst => "0",
      q(0) => register9_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x68,
      clk => clk_1_sg_x68,
      d => register8_q_net,
      en => "1",
      rst(0) => inverter1_op_net,
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/End of Tx Ctrl"

entity end_of_tx_ctrl_entity_87a363d0f3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fifo_emtpy: in std_logic; 
    tx_reset: in std_logic; 
    tx_started: in std_logic; 
    output_en: out std_logic
  );
end end_of_tx_ctrl_entity_87a363d0f3;

architecture structural of end_of_tx_ctrl_entity_87a363d0f3 is
  signal ce_1_sg_x72: std_logic;
  signal clk_1_sg_x72: std_logic;
  signal delay2_q_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical_y_net_x34: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x3: std_logic;
  signal relational1_op_net_x1: std_logic;

begin
  ce_1_sg_x72 <= ce_1;
  clk_1_sg_x72 <= clk_1;
  relational1_op_net_x1 <= fifo_emtpy;
  logical_y_net_x34 <= tx_reset;
  register2_q_net_x1 <= tx_started;
  output_en <= register2_q_net_x3;

  delay2: entity work.xldelay
    generic map (
      latency => 4,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x72,
      clk => clk_1_sg_x72,
      d(0) => logical1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net,
      d1(0) => logical_y_net_x34,
      y(0) => logical3_y_net_x0
    );

  posedge1_496317b7f8: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x72,
      clk_1 => clk_1_sg_x72,
      d => relational1_op_net_x1,
      q => logical1_y_net_x0
    );

  posedge_50c201ff09: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x72,
      clk_1 => clk_1_sg_x72,
      d => register2_q_net_x1,
      q => logical1_y_net_x1
    );

  s_r_latch_9b4b04babf: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x72,
      clk_1 => clk_1_sg_x72,
      r => logical3_y_net_x0,
      s => logical1_y_net_x1,
      q => register2_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/FIFO/I/Q Concat"

entity q_concat_entity_9872452a0b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    q: in std_logic_vector(15 downto 0); 
    iq: out std_logic_vector(31 downto 0)
  );
end q_concat_entity_9872452a0b;

architecture structural of q_concat_entity_9872452a0b is
  signal ce_1_sg_x73: std_logic;
  signal clk_1_sg_x73: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert1_dout_net: std_logic_vector(15 downto 0);
  signal convert_dout_net: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x4: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x73 <= ce_1;
  clk_1_sg_x73 <= clk_1;
  reinterpret2_output_port_net_x4 <= i;
  reinterpret3_output_port_net_x4 <= q;
  iq <= concat_y_net_x0;

  concat: entity work.concat_a369e00c6b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net_x0
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x73,
      clk => clk_1_sg_x73,
      clr => '0',
      din => reinterpret2_output_port_net_x4,
      en => "1",
      dout => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x73,
      clk => clk_1_sg_x73,
      clr => '0',
      din => reinterpret3_output_port_net_x4,
      en => "1",
      dout => convert1_dout_net
    );

  reinterpret: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_dout_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert1_dout_net,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/FIFO"

entity fifo_entity_ed2bc31ace is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_i: in std_logic_vector(15 downto 0); 
    fft_q: in std_logic_vector(15 downto 0); 
    rd: in std_logic; 
    reset: in std_logic; 
    tx_reset: in std_logic; 
    write: in std_logic; 
    empty: out std_logic; 
    i: out std_logic_vector(15 downto 0); 
    output_fifo_occ: out std_logic_vector(7 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end fifo_entity_ed2bc31ace;

architecture structural of fifo_entity_ed2bc31ace is
  signal ce_1_sg_x74: std_logic;
  signal clk_1_sg_x74: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant2_op_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal delay1_q_net: std_logic;
  signal delay3_q_net_x2: std_logic;
  signal fifo_dcount_net_x1: std_logic_vector(7 downto 0);
  signal fifo_dout_net_x0: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical4_y_net: std_logic;
  signal logical_y_net_x35: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net_x0: std_logic;
  signal register_q_net: std_logic_vector(31 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x5: std_logic_vector(15 downto 0);
  signal relational1_op_net_x2: std_logic;

begin
  ce_1_sg_x74 <= ce_1;
  clk_1_sg_x74 <= clk_1;
  reinterpret2_output_port_net_x5 <= fft_i;
  reinterpret3_output_port_net_x5 <= fft_q;
  register3_q_net_x0 <= rd;
  logical1_y_net_x0 <= reset;
  logical_y_net_x35 <= tx_reset;
  delay3_q_net_x2 <= write;
  empty <= relational1_op_net_x2;
  i <= reinterpret2_output_port_net_x1;
  output_fifo_occ <= fifo_dcount_net_x1;
  q <= reinterpret3_output_port_net_x1;

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      clr => '0',
      din(0) => logical1_y_net_x0,
      en => "1",
      dout(0) => convert2_dout_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 12,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      d(0) => logical_y_net_x35,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  fifo: entity work.xlfifogen_wlan_phy_tx_pmd
    generic map (
      core_name0 => "fifo_fg92_6a1156e8dc43a711",
      data_count_width => 8,
      data_width => 32,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      din => register_q_net,
      en => '1',
      re => register3_q_net_x0,
      re_ce => ce_1_sg_x74,
      rst => register2_q_net,
      we => register1_q_net,
      we_ce => ce_1_sg_x74,
      dcount => fifo_dcount_net_x1,
      dout => fifo_dout_net_x0
    );

  logical4: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay1_q_net,
      d1(0) => convert2_dout_net,
      y(0) => logical4_y_net
    );

  q_concat_9872452a0b: entity work.q_concat_entity_9872452a0b
    port map (
      ce_1 => ce_1_sg_x74,
      clk_1 => clk_1_sg_x74,
      i => reinterpret2_output_port_net_x5,
      q => reinterpret3_output_port_net_x5,
      iq => concat_y_net_x0
    );

  q_slice_a49b8b75e5: entity work.q_slice_entity_6da961fd0c
    port map (
      iq => fifo_dout_net_x0,
      i => reinterpret2_output_port_net_x1,
      q => reinterpret3_output_port_net_x1
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      d(0) => delay3_q_net_x2,
      en => "1",
      rst => "0",
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      d(0) => logical4_y_net,
      en => "1",
      rst => "0",
      q(0) => register2_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 32,
      init_value => b"00000000000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      d => concat_y_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net
    );

  relational1: entity work.relational_6dad3a03fc
    port map (
      a => fifo_dcount_net_x1,
      b(0) => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/Preamble Gen"

entity preamble_gen_entity_c25e867a97 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    rd_en: in std_logic; 
    tx_reset: in std_logic; 
    tx_running: in std_logic; 
    done: out std_logic; 
    early_done: out std_logic; 
    i: out std_logic_vector(15 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end preamble_gen_entity_c25e867a97;

architecture structural of preamble_gen_entity_c25e867a97 is
  signal ce_1_sg_x76: std_logic;
  signal clk_1_sg_x76: std_logic;
  signal constant3_op_net: std_logic_vector(8 downto 0);
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay4_q_net: std_logic;
  signal inverter1_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical_y_net_x36: std_logic;
  signal preamble_i_data_net: std_logic_vector(15 downto 0);
  signal preamble_q_data_net: std_logic_vector(15 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register2_q_net_x2: std_logic;
  signal register2_q_net_x3: std_logic;
  signal register2_q_net_x4: std_logic_vector(15 downto 0);
  signal register3_q_net_x0: std_logic_vector(15 downto 0);
  signal register_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;

begin
  ce_1_sg_x76 <= ce_1;
  clk_1_sg_x76 <= clk_1;
  register2_q_net_x2 <= rd_en;
  logical_y_net_x36 <= tx_reset;
  register2_q_net_x3 <= tx_running;
  done <= register1_q_net_x0;
  early_done <= register_q_net_x0;
  i <= register2_q_net_x4;
  q <= register3_q_net_x0;

  constant3: entity work.constant_0512fd5e4c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_36e2bb554c95560d",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => delay4_q_net,
      op => counter_op_net
    );

  delay4: entity work.xldelay
    generic map (
      latency => 4,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d(0) => logical_y_net_x36,
      en => '1',
      rst => '1',
      q(0) => delay4_q_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      ip(0) => relational2_op_net,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x3,
      d1(0) => register2_q_net_x2,
      d2(0) => relational2_op_net,
      y(0) => logical1_y_net
    );

  preamble_i: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 9,
      c_address_width => 9,
      c_width => 16,
      core_name0 => "dmg_72_d16d082a6bc00ceb",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      en => "1",
      data => preamble_i_data_net
    );

  preamble_q: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 9,
      c_address_width => 9,
      c_width => 16,
      core_name0 => "dmg_72_2b0650236539a42c",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      en => "1",
      data => preamble_q_data_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d(0) => register_q_net_x0,
      en(0) => register2_q_net_x2,
      rst(0) => delay4_q_net,
      q(0) => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d => preamble_i_data_net,
      en(0) => register2_q_net_x2,
      rst(0) => delay4_q_net,
      q => register2_q_net_x4
    );

  register3: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d => preamble_q_data_net,
      en(0) => register2_q_net_x2,
      rst(0) => delay4_q_net,
      q => register3_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d(0) => inverter1_op_net,
      en(0) => register2_q_net_x2,
      rst(0) => delay4_q_net,
      q(0) => register_q_net_x0
    );

  relational2: entity work.relational_82fb466a8b
    port map (
      a => counter_op_net,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/Scaling"

entity scaling_entity_a269710a35 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    payload_i: in std_logic_vector(15 downto 0); 
    payload_q: in std_logic_vector(15 downto 0); 
    payload_sel: in std_logic; 
    preamble_i: in std_logic_vector(15 downto 0); 
    preamble_q: in std_logic_vector(15 downto 0); 
    regtx_scaling_payload: in std_logic_vector(15 downto 0); 
    regtx_scaling_preamble: in std_logic_vector(15 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end scaling_entity_a269710a35;

architecture structural of scaling_entity_a269710a35 is
  signal ce_1_sg_x78: std_logic;
  signal clk_1_sg_x78: std_logic;
  signal mult1_p_net_x1: std_logic_vector(11 downto 0);
  signal mult_p_net_x1: std_logic_vector(11 downto 0);
  signal mux1_y_net: std_logic_vector(15 downto 0);
  signal mux2_y_net: std_logic_vector(15 downto 0);
  signal mux_y_net: std_logic_vector(15 downto 0);
  signal register13_q_net_x0: std_logic_vector(15 downto 0);
  signal register14_q_net_x0: std_logic_vector(15 downto 0);
  signal register1_q_net: std_logic_vector(15 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register2_q_net_x5: std_logic_vector(15 downto 0);
  signal register3_q_net_x1: std_logic_vector(15 downto 0);
  signal register5_q_net: std_logic;
  signal register8_q_net: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x78 <= ce_1;
  clk_1_sg_x78 <= clk_1;
  reinterpret2_output_port_net_x2 <= payload_i;
  reinterpret3_output_port_net_x2 <= payload_q;
  register1_q_net_x1 <= payload_sel;
  register2_q_net_x5 <= preamble_i;
  register3_q_net_x1 <= preamble_q;
  register14_q_net_x0 <= regtx_scaling_payload;
  register13_q_net_x0 <= regtx_scaling_preamble;
  i <= mult_p_net_x1;
  q <= mult1_p_net_x1;

  mult: entity work.xlmult_wlan_phy_tx_pmd
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 15,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 12,
      b_width => 16,
      c_a_type => 0,
      c_a_width => 16,
      c_b_type => 1,
      c_b_width => 16,
      c_baat => 16,
      c_output_width => 32,
      c_type => 0,
      core_name0 => "mult_11_2_f2bb5a57782af7d9",
      extra_registers => 1,
      multsign => 2,
      overflow => 2,
      p_arith => xlSigned,
      p_bin_pt => 11,
      p_width => 12,
      quantization => 1
    )
    port map (
      a => register8_q_net,
      b => mux1_y_net,
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      core_ce => ce_1_sg_x78,
      core_clk => clk_1_sg_x78,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult_p_net_x1
    );

  mult1: entity work.xlmult_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 12,
      a_width => 16,
      b_arith => xlSigned,
      b_bin_pt => 15,
      b_width => 16,
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 0,
      c_b_width => 16,
      c_baat => 16,
      c_output_width => 32,
      c_type => 0,
      core_name0 => "mult_11_2_414c0fa5acc33f35",
      extra_registers => 1,
      multsign => 2,
      overflow => 2,
      p_arith => xlSigned,
      p_bin_pt => 11,
      p_width => 12,
      quantization => 1
    )
    port map (
      a => mux1_y_net,
      b => register1_q_net,
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      core_ce => ce_1_sg_x78,
      core_clk => clk_1_sg_x78,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult1_p_net_x1
    );

  mux: entity work.mux_a54904b290
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register2_q_net_x5,
      d1 => reinterpret2_output_port_net_x2,
      sel(0) => register1_q_net_x1,
      y => mux_y_net
    );

  mux1: entity work.mux_a54904b290
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register14_q_net_x0,
      d1 => register13_q_net_x0,
      sel(0) => register5_q_net,
      y => mux1_y_net
    );

  mux2: entity work.mux_a54904b290
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register3_q_net_x1,
      d1 => reinterpret3_output_port_net_x2,
      sel(0) => register1_q_net_x1,
      y => mux2_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      d => mux2_y_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      d(0) => register1_q_net_x1,
      en => "1",
      rst => "0",
      q(0) => register5_q_net
    );

  register8: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      d => mux_y_net,
      en => "1",
      rst => "0",
      q => register8_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs"

entity \preamble___outputs_entity_82fcc722dc\ is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    iq_tvalid: in std_logic; 
    q: in std_logic_vector(15 downto 0); 
    register1: in std_logic_vector(3 downto 0); 
    register13: in std_logic_vector(15 downto 0); 
    register14: in std_logic_vector(15 downto 0); 
    register23: in std_logic; 
    register3_x0: in std_logic; 
    register4_x0: in std_logic; 
    register5: in std_logic; 
    register6: in std_logic; 
    tx_iq_samp_ce: in std_logic; 
    tx_reset: in std_logic; 
    tx_start: in std_logic; 
    dac_outputs: out std_logic_vector(11 downto 0); 
    dac_outputs_x0: out std_logic_vector(11 downto 0); 
    dac_outputs_x1: out std_logic_vector(11 downto 0); 
    dac_outputs_x2: out std_logic_vector(11 downto 0); 
    dac_outputs_x3: out std_logic_vector(11 downto 0); 
    dac_outputs_x4: out std_logic_vector(11 downto 0); 
    dac_outputs_x5: out std_logic_vector(11 downto 0); 
    dac_outputs_x6: out std_logic_vector(11 downto 0); 
    fifo: out std_logic_vector(7 downto 0); 
    last_samp_output_to_dacs: out std_logic
  );
end \preamble___outputs_entity_82fcc722dc\;

architecture structural of \preamble___outputs_entity_82fcc722dc\ is
  signal ce_1_sg_x79: std_logic;
  signal clk_1_sg_x79: std_logic;
  signal convert2_dout_net_x2: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay3_q_net_x3: std_logic;
  signal fifo_dcount_net_x2: std_logic_vector(7 downto 0);
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical_y_net_x38: std_logic;
  signal mult1_p_net_x1: std_logic_vector(11 downto 0);
  signal mult_p_net_x1: std_logic_vector(11 downto 0);
  signal register13_q_net_x1: std_logic_vector(15 downto 0);
  signal register14_q_net_x1: std_logic_vector(15 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register1_q_net_x4: std_logic_vector(3 downto 0);
  signal register1_q_net_x5: std_logic_vector(11 downto 0);
  signal register23_q_net_x2: std_logic;
  signal register2_q_net_x3: std_logic;
  signal register2_q_net_x4: std_logic;
  signal register2_q_net_x5: std_logic_vector(15 downto 0);
  signal register2_q_net_x6: std_logic;
  signal register2_q_net_x7: std_logic_vector(11 downto 0);
  signal register3_q_net_x0: std_logic;
  signal register3_q_net_x1: std_logic_vector(15 downto 0);
  signal register3_q_net_x5: std_logic;
  signal register3_q_net_x6: std_logic;
  signal register3_q_net_x7: std_logic_vector(11 downto 0);
  signal register4_q_net: std_logic;
  signal register4_q_net_x3: std_logic;
  signal register4_q_net_x4: std_logic_vector(11 downto 0);
  signal register5_q_net_x3: std_logic;
  signal register5_q_net_x4: std_logic_vector(11 downto 0);
  signal register6_q_net_x3: std_logic;
  signal register6_q_net_x4: std_logic_vector(11 downto 0);
  signal register7_q_net_x1: std_logic_vector(11 downto 0);
  signal register_q_net_x1: std_logic;
  signal register_q_net_x2: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x6: std_logic_vector(15 downto 0);
  signal relational1_op_net_x2: std_logic;

begin
  ce_1_sg_x79 <= ce_1;
  clk_1_sg_x79 <= clk_1;
  reinterpret2_output_port_net_x6 <= i;
  delay3_q_net_x3 <= iq_tvalid;
  reinterpret3_output_port_net_x6 <= q;
  register1_q_net_x4 <= register1;
  register13_q_net_x1 <= register13;
  register14_q_net_x1 <= register14;
  register23_q_net_x2 <= register23;
  register3_q_net_x5 <= register3_x0;
  register4_q_net_x3 <= register4_x0;
  register5_q_net_x3 <= register5;
  register6_q_net_x3 <= register6;
  convert2_dout_net_x2 <= tx_iq_samp_ce;
  logical_y_net_x38 <= tx_reset;
  register3_q_net_x6 <= tx_start;
  dac_outputs <= register_q_net_x2;
  dac_outputs_x0 <= register1_q_net_x5;
  dac_outputs_x1 <= register2_q_net_x7;
  dac_outputs_x2 <= register3_q_net_x7;
  dac_outputs_x3 <= register4_q_net_x4;
  dac_outputs_x4 <= register5_q_net_x4;
  dac_outputs_x5 <= register6_q_net_x4;
  dac_outputs_x6 <= register7_q_net_x1;
  fifo <= fifo_dcount_net_x2;
  last_samp_output_to_dacs <= delay2_q_net_x0;

  dac_outputs_fec48642b9: entity work.dac_outputs_entity_fec48642b9
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      en => register2_q_net_x3,
      i => mult_p_net_x1,
      q => mult1_p_net_x1,
      register1_x0 => register1_q_net_x4,
      register23 => register23_q_net_x2,
      register3_x0 => register3_q_net_x5,
      register4_x0 => register4_q_net_x3,
      register5_x0 => register5_q_net_x3,
      register6_x0 => register6_q_net_x3,
      register1_x1 => register1_q_net_x5,
      register2_x0 => register2_q_net_x7,
      register3_x1 => register3_q_net_x7,
      register4_x1 => register4_q_net_x4,
      register5_x1 => register5_q_net_x4,
      register6_x1 => register6_q_net_x4,
      register7_x0 => register7_q_net_x1,
      register_x1 => register_q_net_x2
    );

  delay2: entity work.xldelay
    generic map (
      latency => 12,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => logical3_y_net,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  end_of_tx_ctrl_87a363d0f3: entity work.end_of_tx_ctrl_entity_87a363d0f3
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      fifo_emtpy => relational1_op_net_x2,
      tx_reset => logical_y_net_x38,
      tx_started => register2_q_net_x4,
      output_en => register2_q_net_x3
    );

  fifo_ed2bc31ace: entity work.fifo_entity_ed2bc31ace
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      fft_i => reinterpret2_output_port_net_x6,
      fft_q => reinterpret3_output_port_net_x6,
      rd => register3_q_net_x0,
      reset => logical1_y_net_x2,
      tx_reset => logical_y_net_x38,
      write => delay3_q_net_x3,
      empty => relational1_op_net_x2,
      i => reinterpret2_output_port_net_x2,
      output_fifo_occ => fifo_dcount_net_x2,
      q => reinterpret3_output_port_net_x2
    );

  logical2: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register_q_net_x1,
      d1(0) => register2_q_net_x4,
      d2(0) => convert2_dout_net_x2,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x2,
      d1(0) => register4_q_net,
      y(0) => logical3_y_net
    );

  posedge_35705d73cb: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      d => register3_q_net_x6,
      q => logical1_y_net_x2
    );

  preamble_gen_c25e867a97: entity work.preamble_gen_entity_c25e867a97
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      rd_en => register2_q_net_x6,
      tx_reset => logical_y_net_x38,
      tx_running => register2_q_net_x4,
      done => register1_q_net_x1,
      early_done => register_q_net_x1,
      i => register2_q_net_x5,
      q => register3_q_net_x1
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => convert2_dout_net_x2,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x6
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => logical2_y_net,
      en => "1",
      rst => "0",
      q(0) => register3_q_net_x0
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => logical2_y_net,
      en => "1",
      rst => "0",
      q(0) => register4_q_net
    );

  s_r_latch_c320bee3e4: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      r => logical_y_net_x38,
      s => logical1_y_net_x2,
      q => register2_q_net_x4
    );

  scaling_a269710a35: entity work.scaling_entity_a269710a35
    port map (
      ce_1 => ce_1_sg_x79,
      clk_1 => clk_1_sg_x79,
      payload_i => reinterpret2_output_port_net_x2,
      payload_q => reinterpret3_output_port_net_x2,
      payload_sel => register1_q_net_x1,
      preamble_i => register2_q_net_x5,
      preamble_q => register3_q_net_x1,
      regtx_scaling_payload => register14_q_net_x1,
      regtx_scaling_preamble => register13_q_net_x1,
      i => mult_p_net_x1,
      q => mult1_p_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Radio Controller & MAC IO"

entity \radio_controller___mac_io_entity_c70eccdf43\ is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    phy_tx_start: in std_logic; 
    rc_phy_start: in std_logic; 
    mac_io_phy_tx_start: out std_logic; 
    rc_io_phy_start: out std_logic
  );
end \radio_controller___mac_io_entity_c70eccdf43\;

architecture structural of \radio_controller___mac_io_entity_c70eccdf43\ is
  signal ce_1_sg_x80: std_logic;
  signal clk_1_sg_x80: std_logic;
  signal convert1_dout_net_x0: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal phy_tx_start_net_x0: std_logic;
  signal rc_phy_start_net_x0: std_logic;

begin
  ce_1_sg_x80 <= ce_1;
  clk_1_sg_x80 <= clk_1;
  phy_tx_start_net_x0 <= phy_tx_start;
  rc_phy_start_net_x0 <= rc_phy_start;
  mac_io_phy_tx_start <= convert1_dout_net_x0;
  rc_io_phy_start <= convert2_dout_net_x0;

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x80,
      clk => clk_1_sg_x80,
      clr => '0',
      din(0) => phy_tx_start_net_x0,
      en => "1",
      dout(0) => convert1_dout_net_x0
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x80,
      clk => clk_1_sg_x80,
      clr => '0',
      din(0) => rc_phy_start_net_x0,
      en => "1",
      dout(0) => convert2_dout_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Registers/Status Bits"

entity status_bits_entity_a326423b7c is
  port (
    regtx_tx_running: in std_logic; 
    x32b: out std_logic_vector(31 downto 0)
  );
end status_bits_entity_a326423b7c;

architecture structural of status_bits_entity_a326423b7c is
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant_op_net: std_logic_vector(30 downto 0);
  signal register2_q_net_x0: std_logic;

begin
  register2_q_net_x0 <= regtx_tx_running;
  x32b <= concat_y_net_x0;

  concat: entity work.concat_e25f797841
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant_op_net,
      in1(0) => register2_q_net_x0,
      y => concat_y_net_x0
    );

  constant_x0: entity work.constant_bc7a810978
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Registers"

entity registers_entity_2d8965b1e5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    from_register1: in std_logic_vector(31 downto 0); 
    from_register2: in std_logic_vector(31 downto 0); 
    from_register3: in std_logic_vector(31 downto 0); 
    from_register4: in std_logic_vector(31 downto 0); 
    from_register5: in std_logic_vector(31 downto 0); 
    from_register6: in std_logic_vector(31 downto 0); 
    register2_x0: in std_logic; 
    constant_x1: out std_logic; 
    register20_x0: out std_logic_vector(31 downto 0); 
    regtx_anta_tx_en: out std_logic; 
    regtx_antb_tx_en: out std_logic; 
    regtx_antc_tx_en: out std_logic; 
    regtx_antd_tx_en: out std_logic; 
    regtx_cp_len: out std_logic_vector(7 downto 0); 
    regtx_fft_scaling: out std_logic_vector(5 downto 0); 
    regtx_num_sc: out std_logic_vector(7 downto 0); 
    regtx_pkt_buf_addr_offset: out std_logic_vector(7 downto 0); 
    regtx_pkt_buf_sel: out std_logic_vector(3 downto 0); 
    regtx_posttx_extension: out std_logic_vector(9 downto 0); 
    regtx_posttx_rf_en_extension: out std_logic_vector(9 downto 0); 
    regtx_posttx_rxsig_valid: out std_logic_vector(9 downto 0); 
    regtx_rc_rxen_enable: out std_logic; 
    regtx_reset: out std_logic; 
    regtx_reset_scrambling_lfsr_perpkt: out std_logic; 
    regtx_scaling_payload: out std_logic_vector(15 downto 0); 
    regtx_scaling_preamble: out std_logic_vector(15 downto 0); 
    regtx_start_direct: out std_logic; 
    regtx_start_indirect: out std_logic; 
    regtx_sw_tx_phy_mode: out std_logic_vector(2 downto 0); 
    regtx_txrunning_output_sel: out std_logic; 
    regtx_use_mac_ant_masks: out std_logic
  );
end registers_entity_2d8965b1e5;

architecture structural of registers_entity_2d8965b1e5 is
  signal b_0_1_y_net: std_logic;
  signal b_14_12_y_net: std_logic_vector(2 downto 0);
  signal b_15_0_y_net: std_logic_vector(15 downto 0);
  signal b_15_8_y_net: std_logic_vector(7 downto 0);
  signal b_19_10_y_net: std_logic_vector(9 downto 0);
  signal b_1_y_net: std_logic;
  signal b_1_y_net_x0: std_logic;
  signal b_23_16_y_net: std_logic_vector(7 downto 0);
  signal b_29_20_y_net: std_logic_vector(9 downto 0);
  signal b_29_24_y_net: std_logic_vector(5 downto 0);
  signal b_2_y_net: std_logic;
  signal b_31_16_y_net: std_logic_vector(15 downto 0);
  signal b_31_y_net: std_logic;
  signal b_3_0_y_net: std_logic_vector(3 downto 0);
  signal b_3_y_net: std_logic;
  signal b_4_y_net: std_logic;
  signal b_5_y_net: std_logic;
  signal b_6_y_net: std_logic;
  signal b_7_0_y_net: std_logic_vector(7 downto 0);
  signal b_7_y_net: std_logic;
  signal b_9_0_y_net: std_logic_vector(9 downto 0);
  signal ce_1_sg_x81: std_logic;
  signal clk_1_sg_x81: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant_op_net_x0: std_logic;
  signal from_register1_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register2_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register3_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register4_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register5_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register6_data_out_net_x0: std_logic_vector(31 downto 0);
  signal lsb_y_net: std_logic;
  signal register10_q_net_x2: std_logic_vector(5 downto 0);
  signal register11_q_net_x0: std_logic;
  signal register12_q_net_x0: std_logic;
  signal register13_q_net_x2: std_logic_vector(15 downto 0);
  signal register14_q_net_x2: std_logic_vector(15 downto 0);
  signal register15_q_net_x0: std_logic_vector(3 downto 0);
  signal register16_q_net_x3: std_logic_vector(7 downto 0);
  signal register17_q_net_x0: std_logic_vector(9 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register20_q_net_x0: std_logic_vector(31 downto 0);
  signal register23_q_net_x3: std_logic;
  signal register24_q_net_x0: std_logic;
  signal register26_q_net_x0: std_logic_vector(2 downto 0);
  signal register27_q_net_x0: std_logic_vector(9 downto 0);
  signal register28_q_net_x0: std_logic_vector(9 downto 0);
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x6: std_logic;
  signal register3_q_net_x6: std_logic;
  signal register4_q_net_x4: std_logic;
  signal register5_q_net_x4: std_logic;
  signal register6_q_net_x4: std_logic;
  signal register7_q_net_x0: std_logic;
  signal register8_q_net_x9: std_logic_vector(7 downto 0);
  signal register9_q_net_x3: std_logic_vector(7 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x81 <= ce_1;
  clk_1_sg_x81 <= clk_1;
  from_register1_data_out_net_x0 <= from_register1;
  from_register2_data_out_net_x0 <= from_register2;
  from_register3_data_out_net_x0 <= from_register3;
  from_register4_data_out_net_x0 <= from_register4;
  from_register5_data_out_net_x0 <= from_register5;
  from_register6_data_out_net_x0 <= from_register6;
  register2_q_net_x1 <= register2_x0;
  constant_x1 <= constant_op_net_x0;
  register20_x0 <= register20_q_net_x0;
  regtx_anta_tx_en <= register3_q_net_x6;
  regtx_antb_tx_en <= register4_q_net_x4;
  regtx_antc_tx_en <= register5_q_net_x4;
  regtx_antd_tx_en <= register6_q_net_x4;
  regtx_cp_len <= register9_q_net_x3;
  regtx_fft_scaling <= register10_q_net_x2;
  regtx_num_sc <= register8_q_net_x9;
  regtx_pkt_buf_addr_offset <= register16_q_net_x3;
  regtx_pkt_buf_sel <= register15_q_net_x0;
  regtx_posttx_extension <= register17_q_net_x0;
  regtx_posttx_rf_en_extension <= register27_q_net_x0;
  regtx_posttx_rxsig_valid <= register28_q_net_x0;
  regtx_rc_rxen_enable <= register1_q_net_x0;
  regtx_reset <= register7_q_net_x0;
  regtx_reset_scrambling_lfsr_perpkt <= register2_q_net_x6;
  regtx_scaling_payload <= register14_q_net_x2;
  regtx_scaling_preamble <= register13_q_net_x2;
  regtx_start_direct <= register11_q_net_x0;
  regtx_start_indirect <= register12_q_net_x0;
  regtx_sw_tx_phy_mode <= register26_q_net_x0;
  regtx_txrunning_output_sel <= register24_q_net_x0;
  regtx_use_mac_ant_masks <= register23_q_net_x3;

  b_0_1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_0_1_y_net
    );

  b_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_1_y_net
    );

  b_14_12: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 14,
      x_width => 32,
      y_width => 3
    )
    port map (
      x => from_register5_data_out_net_x0,
      y => b_14_12_y_net
    );

  b_15_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 15,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => from_register3_data_out_net_x0,
      y => b_15_0_y_net
    );

  b_15_8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_15_8_y_net
    );

  b_19_10: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 19,
      x_width => 32,
      y_width => 10
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_19_10_y_net
    );

  b_1_x0: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register2_data_out_net_x0,
      y(0) => b_1_y_net_x0
    );

  b_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_2_y_net
    );

  b_23_16: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register4_data_out_net_x0,
      y => b_23_16_y_net
    );

  b_29_20: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 29,
      x_width => 32,
      y_width => 10
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_29_20_y_net
    );

  b_29_24: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 29,
      x_width => 32,
      y_width => 6
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_29_24_y_net
    );

  b_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_3_y_net
    );

  b_31: entity work.xlslice
    generic map (
      new_lsb => 31,
      new_msb => 31,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_31_y_net
    );

  b_31_16: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 31,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => from_register3_data_out_net_x0,
      y => b_31_16_y_net
    );

  b_3_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 32,
      y_width => 4
    )
    port map (
      x => from_register4_data_out_net_x0,
      y => b_3_0_y_net
    );

  b_4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_4_y_net
    );

  b_5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_5_y_net
    );

  b_6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_6_y_net
    );

  b_7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_7_y_net
    );

  b_7_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_7_0_y_net
    );

  b_9_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 32,
      y_width => 10
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_9_0_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net_x0
    );

  lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register2_data_out_net_x0,
      y(0) => lsb_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_0_1_y_net,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register10: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_29_24_y_net,
      en => "1",
      rst => "0",
      q => register10_q_net_x2
    );

  register11: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => lsb_y_net,
      en => "1",
      rst => "0",
      q(0) => register11_q_net_x0
    );

  register12: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_1_y_net_x0,
      en => "1",
      rst => "0",
      q(0) => register12_q_net_x0
    );

  register13: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => reinterpret_output_port_net,
      en => "1",
      rst => "0",
      q => register13_q_net_x2
    );

  register14: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => reinterpret1_output_port_net,
      en => "1",
      rst => "0",
      q => register14_q_net_x2
    );

  register15: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_3_0_y_net,
      en => "1",
      rst => "0",
      q => register15_q_net_x0
    );

  register16: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_23_16_y_net,
      en => "1",
      rst => "0",
      q => register16_q_net_x3
    );

  register17: entity work.xlregister
    generic map (
      d_width => 10,
      init_value => b"0000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_9_0_y_net,
      en => "1",
      rst => "0",
      q => register17_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_1_y_net,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x6
    );

  register20: entity work.xlregister
    generic map (
      d_width => 32,
      init_value => b"00000000000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => concat_y_net_x0,
      en => "1",
      rst => "0",
      q => register20_q_net_x0
    );

  register23: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_6_y_net,
      en => "1",
      rst => "0",
      q(0) => register23_q_net_x3
    );

  register24: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_7_y_net,
      en => "1",
      rst => "0",
      q(0) => register24_q_net_x0
    );

  register26: entity work.xlregister
    generic map (
      d_width => 3,
      init_value => b"000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_14_12_y_net,
      en => "1",
      rst => "0",
      q => register26_q_net_x0
    );

  register27: entity work.xlregister
    generic map (
      d_width => 10,
      init_value => b"0000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_19_10_y_net,
      en => "1",
      rst => "0",
      q => register27_q_net_x0
    );

  register28: entity work.xlregister
    generic map (
      d_width => 10,
      init_value => b"0000000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_29_20_y_net,
      en => "1",
      rst => "0",
      q => register28_q_net_x0
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_2_y_net,
      en => "1",
      rst => "0",
      q(0) => register3_q_net_x6
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_3_y_net,
      en => "1",
      rst => "0",
      q(0) => register4_q_net_x4
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_4_y_net,
      en => "1",
      rst => "0",
      q(0) => register5_q_net_x4
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_5_y_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x4
    );

  register7: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d(0) => b_31_y_net,
      en => "1",
      rst => "0",
      q(0) => register7_q_net_x0
    );

  register8: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_7_0_y_net,
      en => "1",
      rst => "0",
      q => register8_q_net_x9
    );

  register9: entity work.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => b_15_8_y_net,
      en => "1",
      rst => "0",
      q => register9_q_net_x3
    );

  reinterpret: entity work.reinterpret_ddc3ebdd7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => b_15_0_y_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_ddc3ebdd7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => b_31_16_y_net,
      output_port => reinterpret1_output_port_net
    );

  status_bits_a326423b7c: entity work.status_bits_entity_a326423b7c
    port map (
      regtx_tx_running => register2_q_net_x1,
      x32b => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Resets"

entity resets_entity_24d0a1b807 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    last_samp_output_to_dacs: in std_logic; 
    regtx_reset: in std_logic; 
    tx_sig_decode_error: in std_logic; 
    tx_force_reset: out std_logic; 
    tx_phy_done: out std_logic; 
    tx_reset: out std_logic
  );
end resets_entity_24d0a1b807;

architecture structural of resets_entity_24d0a1b807 is
  signal ce_1_sg_x84: std_logic;
  signal clk_1_sg_x84: std_logic;
  signal constant_op_net: std_logic;
  signal convert1_dout_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay_q_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical4_y_net_x9: std_logic;
  signal logical_y_net_x39: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register7_q_net_x1: std_logic;
  signal simulation_multiplexer_dout_net: std_logic;

begin
  ce_1_sg_x84 <= ce_1;
  clk_1_sg_x84 <= clk_1;
  delay2_q_net_x1 <= last_samp_output_to_dacs;
  register7_q_net_x1 <= regtx_reset;
  logical4_y_net_x9 <= tx_sig_decode_error;
  tx_force_reset <= convert1_dout_net_x0;
  tx_phy_done <= logical1_y_net_x4;
  tx_reset <= logical_y_net_x39;

  constant_x0: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x84,
      clk => clk_1_sg_x84,
      clr => '0',
      din(0) => register7_q_net_x1,
      en => "1",
      dout(0) => convert1_dout_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 16,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x84,
      clk => clk_1_sg_x84,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x0
    );

  logical: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => simulation_multiplexer_dout_net,
      d1(0) => convert1_dout_net_x0,
      d2(0) => register2_q_net_x0,
      y(0) => logical_y_net_x39
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net_x1,
      d1(0) => logical4_y_net_x9,
      y(0) => logical1_y_net_x1
    );

  posedge1_cd01046e00: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x84,
      clk_1 => clk_1_sg_x84,
      d => logical1_y_net_x1,
      q => logical1_y_net_x4
    );

  s_r_latch_3226b7fe2e: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x84,
      clk_1 => clk_1_sg_x84,
      r => delay_q_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x0
    );

  simulation_multiplexer: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => constant_op_net,
      dout(0) => simulation_multiplexer_dout_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Sampling Clock"

entity sampling_clock_entity_a1a467035e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    samp_ce: in std_logic; 
    tx_iq_samp_ce: out std_logic
  );
end sampling_clock_entity_a1a467035e;

architecture structural of sampling_clock_entity_a1a467035e is
  signal ce_1_sg_x85: std_logic;
  signal clk_1_sg_x85: std_logic;
  signal convert2_dout_net_x3: std_logic;
  signal samp_ce_net_x0: std_logic;

begin
  ce_1_sg_x85 <= ce_1;
  clk_1_sg_x85 <= clk_1;
  samp_ce_net_x0 <= samp_ce;
  tx_iq_samp_ce <= convert2_dout_net_x3;

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      din(0) => samp_ce_net_x0,
      en => "1",
      dout(0) => convert2_dout_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Add MAC Extension"

entity add_mac_extension_entity_ff6c76ae09 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    iq_done: in std_logic; 
    regtx_posttx_extension: in std_logic_vector(9 downto 0); 
    tx_force_reset: in std_logic; 
    tx_iq_samp_ce: in std_logic; 
    tx_start: in std_logic; 
    tx_active: out std_logic
  );
end add_mac_extension_entity_ff6c76ae09;

architecture structural of add_mac_extension_entity_ff6c76ae09 is
  signal ce_1_sg_x88: std_logic;
  signal clk_1_sg_x88: std_logic;
  signal convert1_dout_net_x1: std_logic;
  signal convert2_dout_net_x4: std_logic;
  signal counter1_op_net: std_logic_vector(9 downto 0);
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal register17_q_net_x1: std_logic_vector(9 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x2: std_logic;
  signal register3_q_net_x8: std_logic;
  signal relational3_op_net: std_logic;

begin
  ce_1_sg_x88 <= ce_1;
  clk_1_sg_x88 <= clk_1;
  logical1_y_net_x6 <= iq_done;
  register17_q_net_x1 <= regtx_posttx_extension;
  convert1_dout_net_x1 <= tx_force_reset;
  convert2_dout_net_x4 <= tx_iq_samp_ce;
  register3_q_net_x8 <= tx_start;
  tx_active <= register2_q_net_x2;

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => logical2_y_net_x1,
      op => counter1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => convert2_dout_net_x4,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => convert1_dout_net_x1,
      y(0) => logical2_y_net_x1
    );

  relational3: entity work.relational_e83dd85005
    port map (
      a => counter1_op_net,
      b => register17_q_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_2da9223410: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      r => logical2_y_net_x1,
      s => logical1_y_net_x6,
      q => register2_q_net_x0
    );

  s_r_latch2_e6ced2723e: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      r => logical2_y_net_x1,
      s => register3_q_net_x8,
      q => register2_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Add TXEN Extension"

entity add_txen_extension_entity_c448d7d5a8 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    iq_done: in std_logic; 
    regtx_posttx_rf_en_extension: in std_logic_vector(9 downto 0); 
    regtx_posttx_rxsig_valid: in std_logic_vector(9 downto 0); 
    tx_force_reset: in std_logic; 
    tx_iq_samp_ce: in std_logic; 
    disable_rf_tx: out std_logic; 
    rxsig_valid: out std_logic
  );
end add_txen_extension_entity_c448d7d5a8;

architecture structural of add_txen_extension_entity_c448d7d5a8 is
  signal ce_1_sg_x93: std_logic;
  signal clk_1_sg_x93: std_logic;
  signal convert1_dout_net_x2: std_logic;
  signal convert2_dout_net_x5: std_logic;
  signal counter1_op_net: std_logic_vector(9 downto 0);
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x10: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x9: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal register27_q_net_x1: std_logic_vector(9 downto 0);
  signal register28_q_net_x1: std_logic_vector(9 downto 0);
  signal register2_q_net_x0: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal relational3_op_net: std_logic;

begin
  ce_1_sg_x93 <= ce_1;
  clk_1_sg_x93 <= clk_1;
  logical1_y_net_x9 <= iq_done;
  register27_q_net_x1 <= regtx_posttx_rf_en_extension;
  register28_q_net_x1 <= regtx_posttx_rxsig_valid;
  convert1_dout_net_x2 <= tx_force_reset;
  convert2_dout_net_x5 <= tx_iq_samp_ce;
  disable_rf_tx <= logical1_y_net_x10;
  rxsig_valid <= logical1_y_net_x11;

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x93,
      clk => clk_1_sg_x93,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => logical2_y_net_x0,
      op => counter1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => convert2_dout_net_x5,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x0,
      d1(0) => convert1_dout_net_x2,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x0,
      d1(0) => relational3_op_net,
      y(0) => logical3_y_net_x0
    );

  posedge1_c7c0a906d1: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x93,
      clk_1 => clk_1_sg_x93,
      d => logical1_y_net_x9,
      q => logical1_y_net_x1
    );

  posedge2_43a5fd301b: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x93,
      clk_1 => clk_1_sg_x93,
      d => logical3_y_net_x0,
      q => logical1_y_net_x10
    );

  posedge3_cf2f9857fd: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x93,
      clk_1 => clk_1_sg_x93,
      d => relational1_op_net_x0,
      q => logical1_y_net_x11
    );

  relational1: entity work.relational_e83dd85005
    port map (
      a => counter1_op_net,
      b => register28_q_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  relational3: entity work.relational_e83dd85005
    port map (
      a => counter1_op_net,
      b => register27_q_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_41b2f20ce9: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x93,
      clk_1 => clk_1_sg_x93,
      r => logical2_y_net_x0,
      s => logical1_y_net_x1,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/PHY Mode Sel"

entity phy_mode_sel_entity_28481ebfc8 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    hw_tx: in std_logic; 
    mac_io_phy_tx_phy_mode: in std_logic_vector(2 downto 0); 
    regtx_sw_tx_phy_mode: in std_logic_vector(2 downto 0); 
    sw_tx: in std_logic; 
    phy_mode: out std_logic_vector(2 downto 0)
  );
end phy_mode_sel_entity_28481ebfc8;

architecture structural of phy_mode_sel_entity_28481ebfc8 is
  signal ce_1_sg_x94: std_logic;
  signal clk_1_sg_x94: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert1_dout_net_x1: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal mux_y_net_x0: std_logic_vector(2 downto 0);
  signal phy_tx_phy_mode_net_x0: std_logic_vector(2 downto 0);
  signal register1_q_net: std_logic_vector(2 downto 0);
  signal register26_q_net_x1: std_logic_vector(2 downto 0);
  signal register2_q_net: std_logic_vector(2 downto 0);
  signal register3_q_net: std_logic;

begin
  ce_1_sg_x94 <= ce_1;
  clk_1_sg_x94 <= clk_1;
  convert1_dout_net_x1 <= hw_tx;
  phy_tx_phy_mode_net_x0 <= mac_io_phy_tx_phy_mode;
  register26_q_net_x1 <= regtx_sw_tx_phy_mode;
  logical5_y_net_x0 <= sw_tx;
  phy_mode <= mux_y_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      clr => '0',
      din(0) => logical5_y_net_x0,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      clr => '0',
      din(0) => convert1_dout_net_x1,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert_dout_net,
      d1(0) => convert1_dout_net,
      y(0) => logical1_y_net
    );

  mux: entity work.mux_1d1da8e0e2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register1_q_net,
      d1 => register2_q_net,
      sel(0) => register3_q_net,
      y => mux_y_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 3,
      init_value => b"000"
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      d => register26_q_net_x1,
      en(0) => convert_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 3,
      init_value => b"000"
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      d => phy_tx_phy_mode_net_x0,
      en(0) => convert1_dout_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      d(0) => convert1_dout_net,
      en(0) => logical1_y_net,
      rst => "0",
      q(0) => register3_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Pkt Buf Sel"

entity pkt_buf_sel_entity_412d479839 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    hw_tx: in std_logic; 
    mac_io_phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    regtx_pkt_buf_sel: in std_logic_vector(3 downto 0); 
    sw_tx: in std_logic; 
    pkt_buf: out std_logic_vector(3 downto 0)
  );
end pkt_buf_sel_entity_412d479839;

architecture structural of pkt_buf_sel_entity_412d479839 is
  signal ce_1_sg_x95: std_logic;
  signal clk_1_sg_x95: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert1_dout_net_x2: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical5_y_net_x1: std_logic;
  signal mux_y_net_x13: std_logic_vector(3 downto 0);
  signal phy_tx_pkt_buf_net_x0: std_logic_vector(3 downto 0);
  signal register15_q_net_x1: std_logic_vector(3 downto 0);
  signal register1_q_net: std_logic_vector(3 downto 0);
  signal register2_q_net: std_logic_vector(3 downto 0);
  signal register3_q_net: std_logic;

begin
  ce_1_sg_x95 <= ce_1;
  clk_1_sg_x95 <= clk_1;
  convert1_dout_net_x2 <= hw_tx;
  phy_tx_pkt_buf_net_x0 <= mac_io_phy_tx_pkt_buf;
  register15_q_net_x1 <= regtx_pkt_buf_sel;
  logical5_y_net_x1 <= sw_tx;
  pkt_buf <= mux_y_net_x13;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      clr => '0',
      din(0) => logical5_y_net_x1,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      clr => '0',
      din(0) => convert1_dout_net_x2,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert_dout_net,
      d1(0) => convert1_dout_net,
      y(0) => logical1_y_net
    );

  mux: entity work.mux_f9c0f11a18
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register1_q_net,
      d1 => register2_q_net,
      sel(0) => register3_q_net,
      y => mux_y_net_x13
    );

  register1: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      d => register15_q_net_x1,
      en(0) => convert_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      d => phy_tx_pkt_buf_net_x0,
      en(0) => convert1_dout_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      d(0) => convert1_dout_net,
      en(0) => logical1_y_net,
      rst => "0",
      q(0) => register3_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Radio TXEN/RXEN Control"

entity rxen_control_entity_677408d8f6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    mac_tx_ant_mask: in std_logic_vector(3 downto 0); 
    regtx_rc_rxen_enable: in std_logic; 
    regtx_use_mac_ant_masks: in std_logic; 
    rx: in std_logic; 
    tx: in std_logic; 
    rc_io_rxen: out std_logic; 
    rc_io_txen_a: out std_logic; 
    rc_io_txen_b: out std_logic; 
    rc_io_txen_c: out std_logic; 
    rc_io_txen_d: out std_logic
  );
end rxen_control_entity_677408d8f6;

architecture structural of rxen_control_entity_677408d8f6 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal ce_1_sg_x100: std_logic;
  signal clk_1_sg_x100: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert7_dout_net: std_logic;
  signal convert8_dout_net: std_logic;
  signal delay1_q_net: std_logic;
  signal delay_q_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical10_y_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;
  signal logical5_y_net: std_logic;
  signal logical6_y_net: std_logic;
  signal logical7_y_net: std_logic;
  signal logical8_y_net: std_logic;
  signal logical9_y_net: std_logic;
  signal rc_rxen_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register1_q_net_x5: std_logic;
  signal register1_q_net_x6: std_logic_vector(3 downto 0);
  signal register23_q_net_x4: std_logic;
  signal register2_q_net_x2: std_logic;
  signal register2_q_net_x3: std_logic;
  signal register2_q_net_x4: std_logic;
  signal register3_q_net_x0: std_logic;
  signal register5_q_net_x0: std_logic;

begin
  ce_1_sg_x100 <= ce_1;
  clk_1_sg_x100 <= clk_1;
  register1_q_net_x6 <= mac_tx_ant_mask;
  register1_q_net_x5 <= regtx_rc_rxen_enable;
  register23_q_net_x4 <= regtx_use_mac_ant_masks;
  register2_q_net_x3 <= rx;
  register2_q_net_x2 <= tx;
  rc_io_rxen <= rc_rxen_x0;
  rc_io_txen_a <= register5_q_net_x0;
  rc_io_txen_b <= register1_q_net_x0;
  rc_io_txen_c <= register2_q_net_x4;
  rc_io_txen_d <= register3_q_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x6,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x6,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x6,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => register1_q_net_x6,
      y(0) => b3_y_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      din(0) => inverter_op_net,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert7: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      din(0) => logical2_y_net,
      en => "1",
      dout(0) => convert7_dout_net
    );

  convert8: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      din(0) => logical3_y_net,
      en => "1",
      dout(0) => convert8_dout_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 32,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical2_y_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 32,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical3_y_net,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      ip(0) => register23_q_net_x4,
      op(0) => inverter_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      ip(0) => delay_q_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      ip(0) => delay1_q_net,
      op(0) => inverter3_op_net
    );

  logical1: entity work.logical_3e1f051fb7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => b1_y_net,
      y(0) => logical1_y_net
    );

  logical10: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert8_dout_net,
      d1(0) => logical4_y_net,
      y(0) => logical10_y_net
    );

  logical2: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register1_q_net_x5,
      d1(0) => register2_q_net_x3,
      d2(0) => inverter3_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter2_op_net,
      d1(0) => register2_q_net_x2,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_3e1f051fb7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => b0_y_net,
      y(0) => logical4_y_net
    );

  logical5: entity work.logical_3e1f051fb7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => b2_y_net,
      y(0) => logical5_y_net
    );

  logical6: entity work.logical_3e1f051fb7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => b3_y_net,
      y(0) => logical6_y_net
    );

  logical7: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert8_dout_net,
      d1(0) => logical1_y_net,
      y(0) => logical7_y_net
    );

  logical8: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert8_dout_net,
      d1(0) => logical5_y_net,
      y(0) => logical8_y_net
    );

  logical9: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert8_dout_net,
      d1(0) => logical6_y_net,
      y(0) => logical9_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical7_y_net,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical8_y_net,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x4
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical9_y_net,
      en => "1",
      rst => "0",
      q(0) => register3_q_net_x0
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => convert7_dout_net,
      en => "1",
      rst => "0",
      q(0) => rc_rxen_x0
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      d(0) => logical10_y_net,
      en => "1",
      rst => "0",
      q(0) => register5_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/S-R Latch2"

entity s_r_latch2_entity_c31d9fc389 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    r: in std_logic; 
    s: in std_logic; 
    q: out std_logic
  );
end s_r_latch2_entity_c31d9fc389;

architecture structural of s_r_latch2_entity_c31d9fc389 is
  signal ce_1_sg_x103: std_logic;
  signal clk_1_sg_x103: std_logic;
  signal constant1_op_net: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;

begin
  ce_1_sg_x103 <= ce_1;
  clk_1_sg_x103 <= clk_1;
  logical8_y_net_x0 <= r;
  logical1_y_net_x4 <= s;
  q <= register2_q_net_x0;

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x103,
      clk => clk_1_sg_x103,
      clr => '0',
      din(0) => logical8_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x103,
      clk => clk_1_sg_x103,
      clr => '0',
      din(0) => logical1_y_net_x4,
      en => "1",
      dout(0) => convert2_dout_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x103,
      clk => clk_1_sg_x103,
      d(0) => constant1_op_net,
      en(0) => convert2_dout_net,
      rst(0) => convert1_dout_net,
      q(0) => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Tx Active Debug Signal/Dly"

entity dly_entity_5c595a7607 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end dly_entity_5c595a7607;

architecture structural of dly_entity_5c595a7607 is
  signal ce_1_sg_x106: std_logic;
  signal clk_1_sg_x106: std_logic;
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant_op_net: std_logic_vector(15 downto 0);
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal convert_dout_net: std_logic;
  signal counter1_op_net: std_logic_vector(4 downto 0);
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register5_q_net_x1: std_logic;
  signal relational1_op_net_x1: std_logic;
  signal relational_op_net_x0: std_logic;

begin
  ce_1_sg_x106 <= ce_1;
  clk_1_sg_x106 <= clk_1;
  register5_q_net_x1 <= d;
  q <= convert2_dout_net_x0;

  constant1: entity work.constant_1e3d9a52c0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant_x0: entity work.constant_18f2e784b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      din(0) => register2_q_net_x0,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      din(0) => register2_q_net_x1,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      din(0) => register2_q_net_x0,
      en => "1",
      dout(0) => convert2_dout_net_x0
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_511eb7a1af6f3f2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      en(0) => convert1_dout_net,
      rst(0) => relational1_op_net_x1,
      op => counter_op_net
    );

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_87d991c7bcfe987f",
      op_arith => xlUnsigned,
      op_width => 5
    )
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      en(0) => convert_dout_net,
      rst(0) => relational1_op_net_x1,
      op => counter1_op_net
    );

  relational: entity work.relational_e55f8c5d80
    port map (
      a => counter_op_net,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net_x0
    );

  relational1: entity work.relational_60871c3374
    port map (
      a => counter1_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x1
    );

  s_r_latch1_8557c9eefb: entity work.s_r_latch2_entity_c31d9fc389
    port map (
      ce_1 => ce_1_sg_x106,
      clk_1 => clk_1_sg_x106,
      r => relational1_op_net_x1,
      s => relational_op_net_x0,
      q => register2_q_net_x0
    );

  s_r_latch2_a2598f1e39: entity work.s_r_latch2_entity_c31d9fc389
    port map (
      ce_1 => ce_1_sg_x106,
      clk_1 => clk_1_sg_x106,
      r => relational1_op_net_x1,
      s => register5_q_net_x1,
      q => register2_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Tx Active Debug Signal"

entity tx_active_debug_signal_entity_fb88e0bcc4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    regtx_txrunning_output_sel: in std_logic; 
    tx_active: in std_logic; 
    register1_x0: out std_logic
  );
end tx_active_debug_signal_entity_fb88e0bcc4;

architecture structural of tx_active_debug_signal_entity_fb88e0bcc4 is
  signal ce_1_sg_x107: std_logic;
  signal clk_1_sg_x107: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal convert9_dout_net: std_logic;
  signal mux_y_net: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register24_q_net_x1: std_logic;
  signal register2_q_net_x4: std_logic;
  signal register5_q_net_x1: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x107 <= ce_1;
  clk_1_sg_x107 <= clk_1;
  register24_q_net_x1 <= regtx_txrunning_output_sel;
  register2_q_net_x4 <= tx_active;
  register1_x0 <= register1_q_net_x0;

  convert9: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x107,
      clk => clk_1_sg_x107,
      clr => '0',
      din(0) => register5_q_net_x1,
      en => "1",
      dout(0) => convert9_dout_net
    );

  dly_5c595a7607: entity work.dly_entity_5c595a7607
    port map (
      ce_1 => ce_1_sg_x107,
      clk_1 => clk_1_sg_x107,
      d => register5_q_net_x1,
      q => convert2_dout_net_x0
    );

  mux: entity work.mux_112ed141f4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert9_dout_net,
      d1(0) => convert2_dout_net_x0,
      sel(0) => register24_q_net_x1,
      y(0) => mux_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x107,
      clk => clk_1_sg_x107,
      d(0) => register_q_net,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x107,
      clk => clk_1_sg_x107,
      d(0) => register2_q_net_x4,
      en => "1",
      rst => "0",
      q(0) => register5_q_net_x1
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x107,
      clk => clk_1_sg_x107,
      d(0) => mux_y_net,
      en => "1",
      rst => "0",
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Tx Gain"

entity tx_gain_entity_164a39bf58 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    hw_tx: in std_logic; 
    phy_tx_gain_a: in std_logic_vector(5 downto 0); 
    phy_tx_gain_b: in std_logic_vector(5 downto 0); 
    phy_tx_gain_c: in std_logic_vector(5 downto 0); 
    phy_tx_gain_d: in std_logic_vector(5 downto 0); 
    sw_tx: in std_logic; 
    tx_gain_a: out std_logic_vector(5 downto 0); 
    tx_gain_b: out std_logic_vector(5 downto 0); 
    tx_gain_c: out std_logic_vector(5 downto 0); 
    tx_gain_d: out std_logic_vector(5 downto 0)
  );
end tx_gain_entity_164a39bf58;

architecture structural of tx_gain_entity_164a39bf58 is
  signal ce_1_sg_x108: std_logic;
  signal clk_1_sg_x108: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert1_dout_net_x3: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical5_y_net_x2: std_logic;
  signal phy_tx_gain_a_net_x0: std_logic_vector(5 downto 0);
  signal phy_tx_gain_b_net_x0: std_logic_vector(5 downto 0);
  signal phy_tx_gain_c_net_x0: std_logic_vector(5 downto 0);
  signal phy_tx_gain_d_net_x0: std_logic_vector(5 downto 0);
  signal register1_q_net_x0: std_logic_vector(5 downto 0);
  signal register2_q_net: std_logic_vector(5 downto 0);
  signal register3_q_net_x0: std_logic_vector(5 downto 0);
  signal register4_q_net: std_logic_vector(5 downto 0);
  signal register5_q_net_x0: std_logic_vector(5 downto 0);
  signal register6_q_net: std_logic_vector(5 downto 0);
  signal register7_q_net_x0: std_logic_vector(5 downto 0);
  signal register8_q_net: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x108 <= ce_1;
  clk_1_sg_x108 <= clk_1;
  convert1_dout_net_x3 <= hw_tx;
  phy_tx_gain_a_net_x0 <= phy_tx_gain_a;
  phy_tx_gain_b_net_x0 <= phy_tx_gain_b;
  phy_tx_gain_c_net_x0 <= phy_tx_gain_c;
  phy_tx_gain_d_net_x0 <= phy_tx_gain_d;
  logical5_y_net_x2 <= sw_tx;
  tx_gain_a <= register1_q_net_x0;
  tx_gain_b <= register3_q_net_x0;
  tx_gain_c <= register5_q_net_x0;
  tx_gain_d <= register7_q_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      clr => '0',
      din(0) => logical5_y_net_x2,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      clr => '0',
      din(0) => convert1_dout_net_x3,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert_dout_net,
      d1(0) => convert1_dout_net,
      y(0) => logical1_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => register2_q_net,
      en => "1",
      rst => "0",
      q => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => phy_tx_gain_a_net_x0,
      en(0) => logical1_y_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => register4_q_net,
      en => "1",
      rst => "0",
      q => register3_q_net_x0
    );

  register4: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => phy_tx_gain_b_net_x0,
      en(0) => logical1_y_net,
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => register6_q_net,
      en => "1",
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => phy_tx_gain_c_net_x0,
      en(0) => logical1_y_net,
      rst => "0",
      q => register6_q_net
    );

  register7: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => register8_q_net,
      en => "1",
      rst => "0",
      q => register7_q_net_x0
    );

  register8: entity work.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      d => phy_tx_gain_d_net_x0,
      en(0) => logical1_y_net,
      rst => "0",
      q => register8_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl"

entity start_ctrl_entity_3ba2a032ad is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    mac_io_phy_tx_ant_mask: in std_logic_vector(3 downto 0); 
    mac_io_phy_tx_start: in std_logic; 
    phy_tx_gain_a: in std_logic_vector(5 downto 0); 
    phy_tx_gain_b: in std_logic_vector(5 downto 0); 
    phy_tx_gain_c: in std_logic_vector(5 downto 0); 
    phy_tx_gain_d: in std_logic_vector(5 downto 0); 
    phy_tx_phy_mode: in std_logic_vector(2 downto 0); 
    phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    rc_io_phy_start: in std_logic; 
    registers: in std_logic_vector(3 downto 0); 
    registers_x0: in std_logic_vector(9 downto 0); 
    registers_x1: in std_logic; 
    registers_x2: in std_logic; 
    registers_x3: in std_logic_vector(2 downto 0); 
    registers_x4: in std_logic_vector(9 downto 0); 
    registers_x5: in std_logic_vector(9 downto 0); 
    regtx_rc_rxen_enable: in std_logic; 
    regtx_start_direct: in std_logic; 
    regtx_start_indirect: in std_logic; 
    tx_force_reset: in std_logic; 
    tx_iq_samp_ce: in std_logic; 
    tx_phy_done: in std_logic; 
    mac_io_phy_tx_done: out std_logic; 
    mac_io_phy_tx_started: out std_logic; 
    mac_tx_ant_mask: out std_logic_vector(3 downto 0); 
    phy_start: out std_logic; 
    rc_io_tx_gain_a: out std_logic_vector(5 downto 0); 
    rc_io_tx_gain_b: out std_logic_vector(5 downto 0); 
    rc_io_tx_gain_c: out std_logic_vector(5 downto 0); 
    rc_io_tx_gain_d: out std_logic_vector(5 downto 0); 
    register2_x0: out std_logic; 
    regtx_tx_running: out std_logic; 
    rxen_control: out std_logic; 
    rxen_control_x0: out std_logic; 
    rxen_control_x1: out std_logic; 
    rxen_control_x2: out std_logic; 
    rxen_control_x3: out std_logic; 
    tx_active_debug_signal: out std_logic; 
    tx_phy_mode_11ag: out std_logic; 
    tx_phy_mode_11n: out std_logic; 
    tx_phy_mode_11n_ac: out std_logic; 
    tx_pkt_buf_sel: out std_logic_vector(3 downto 0)
  );
end start_ctrl_entity_3ba2a032ad;

architecture structural of start_ctrl_entity_3ba2a032ad is
  signal ce_1_sg_x110: std_logic;
  signal clk_1_sg_x110: std_logic;
  signal convert1_dout_net_x4: std_logic;
  signal convert1_dout_net_x5: std_logic;
  signal convert2_dout_net_x1: std_logic;
  signal convert2_dout_net_x6: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x12: std_logic;
  signal logical1_y_net_x13: std_logic;
  signal logical1_y_net_x14: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical3_y_net_x7: std_logic;
  signal logical4_y_net_x0: std_logic;
  signal logical5_y_net_x2: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical7_y_net_x0: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x0: std_logic_vector(2 downto 0);
  signal mux_y_net_x14: std_logic_vector(3 downto 0);
  signal phy_tx_ant_mask_net_x0: std_logic_vector(3 downto 0);
  signal phy_tx_gain_a_net_x1: std_logic_vector(5 downto 0);
  signal phy_tx_gain_b_net_x1: std_logic_vector(5 downto 0);
  signal phy_tx_gain_c_net_x1: std_logic_vector(5 downto 0);
  signal phy_tx_gain_d_net_x1: std_logic_vector(5 downto 0);
  signal phy_tx_phy_mode_net_x1: std_logic_vector(2 downto 0);
  signal phy_tx_pkt_buf_net_x1: std_logic_vector(3 downto 0);
  signal rc_rxen_x1: std_logic;
  signal register11_q_net_x1: std_logic;
  signal register12_q_net_x1: std_logic;
  signal register15_q_net_x2: std_logic_vector(3 downto 0);
  signal register17_q_net_x2: std_logic_vector(9 downto 0);
  signal register1_q_net_x10: std_logic;
  signal register1_q_net_x11: std_logic_vector(5 downto 0);
  signal register1_q_net_x7: std_logic;
  signal register1_q_net_x8: std_logic;
  signal register1_q_net_x9: std_logic_vector(3 downto 0);
  signal register23_q_net_x5: std_logic;
  signal register24_q_net_x2: std_logic;
  signal register26_q_net_x2: std_logic_vector(2 downto 0);
  signal register27_q_net_x2: std_logic_vector(9 downto 0);
  signal register28_q_net_x2: std_logic_vector(9 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x5: std_logic;
  signal register2_q_net_x6: std_logic;
  signal register2_q_net_x7: std_logic;
  signal register2_q_net_x8: std_logic;
  signal register2_q_net_x9: std_logic;
  signal register3_q_net_x10: std_logic_vector(5 downto 0);
  signal register3_q_net_x2: std_logic;
  signal register3_q_net_x9: std_logic;
  signal register4_q_net: std_logic_vector(3 downto 0);
  signal register5_q_net_x2: std_logic;
  signal register5_q_net_x3: std_logic_vector(5 downto 0);
  signal register7_q_net_x1: std_logic_vector(5 downto 0);
  signal slice1_y_net_x13: std_logic;
  signal slice2_y_net: std_logic;
  signal slice_y_net_x6: std_logic;

begin
  ce_1_sg_x110 <= ce_1;
  clk_1_sg_x110 <= clk_1;
  phy_tx_ant_mask_net_x0 <= mac_io_phy_tx_ant_mask;
  convert1_dout_net_x4 <= mac_io_phy_tx_start;
  phy_tx_gain_a_net_x1 <= phy_tx_gain_a;
  phy_tx_gain_b_net_x1 <= phy_tx_gain_b;
  phy_tx_gain_c_net_x1 <= phy_tx_gain_c;
  phy_tx_gain_d_net_x1 <= phy_tx_gain_d;
  phy_tx_phy_mode_net_x1 <= phy_tx_phy_mode;
  phy_tx_pkt_buf_net_x1 <= phy_tx_pkt_buf;
  convert2_dout_net_x1 <= rc_io_phy_start;
  register15_q_net_x2 <= registers;
  register17_q_net_x2 <= registers_x0;
  register23_q_net_x5 <= registers_x1;
  register24_q_net_x2 <= registers_x2;
  register26_q_net_x2 <= registers_x3;
  register27_q_net_x2 <= registers_x4;
  register28_q_net_x2 <= registers_x5;
  register1_q_net_x7 <= regtx_rc_rxen_enable;
  register11_q_net_x1 <= regtx_start_direct;
  register12_q_net_x1 <= regtx_start_indirect;
  convert1_dout_net_x5 <= tx_force_reset;
  convert2_dout_net_x6 <= tx_iq_samp_ce;
  logical1_y_net_x13 <= tx_phy_done;
  mac_io_phy_tx_done <= logical1_y_net_x14;
  mac_io_phy_tx_started <= logical1_y_net_x6;
  mac_tx_ant_mask <= register1_q_net_x9;
  phy_start <= register3_q_net_x9;
  rc_io_tx_gain_a <= register1_q_net_x11;
  rc_io_tx_gain_b <= register3_q_net_x10;
  rc_io_tx_gain_c <= register5_q_net_x3;
  rc_io_tx_gain_d <= register7_q_net_x1;
  register2_x0 <= register2_q_net_x8;
  regtx_tx_running <= register2_q_net_x9;
  rxen_control <= register1_q_net_x8;
  rxen_control_x0 <= register2_q_net_x7;
  rxen_control_x1 <= register3_q_net_x2;
  rxen_control_x2 <= rc_rxen_x1;
  rxen_control_x3 <= register5_q_net_x2;
  tx_active_debug_signal <= register1_q_net_x10;
  tx_phy_mode_11ag <= slice_y_net_x6;
  tx_phy_mode_11n <= slice1_y_net_x13;
  tx_phy_mode_11n_ac <= logical3_y_net_x7;
  tx_pkt_buf_sel <= mux_y_net_x14;

  add_mac_extension_ff6c76ae09: entity work.add_mac_extension_entity_ff6c76ae09
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      iq_done => logical1_y_net_x13,
      regtx_posttx_extension => register17_q_net_x2,
      tx_force_reset => convert1_dout_net_x5,
      tx_iq_samp_ce => convert2_dout_net_x6,
      tx_start => register3_q_net_x9,
      tx_active => register2_q_net_x5
    );

  add_txen_extension_c448d7d5a8: entity work.add_txen_extension_entity_c448d7d5a8
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      iq_done => logical1_y_net_x13,
      regtx_posttx_rf_en_extension => register27_q_net_x2,
      regtx_posttx_rxsig_valid => register28_q_net_x2,
      tx_force_reset => convert1_dout_net_x5,
      tx_iq_samp_ce => convert2_dout_net_x6,
      disable_rf_tx => logical1_y_net_x11,
      rxsig_valid => logical1_y_net_x12
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register11_q_net_x1,
      d1(0) => convert2_dout_net_x1,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register12_q_net_x1,
      d1(0) => convert1_dout_net_x4,
      y(0) => logical1_y_net_x1
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => slice1_y_net_x13,
      d1(0) => slice2_y_net,
      y(0) => logical3_y_net_x7
    );

  logical4: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x2,
      d1(0) => logical1_y_net_x3,
      y(0) => logical4_y_net_x0
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register12_q_net_x1,
      d1(0) => register11_q_net_x1,
      y(0) => logical5_y_net_x2
    );

  logical6: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical4_y_net_x0,
      d1(0) => convert1_dout_net_x5,
      y(0) => logical6_y_net_x0
    );

  logical7: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x4,
      d1(0) => convert1_dout_net_x5,
      y(0) => logical7_y_net_x0
    );

  logical8: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x12,
      d1(0) => convert1_dout_net_x5,
      y(0) => logical8_y_net_x0
    );

  negedge_5ee9de3524: entity work.negedge_entity_02af90a306
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      d => register2_q_net_x5,
      q => logical1_y_net_x14
    );

  phy_mode_sel_28481ebfc8: entity work.phy_mode_sel_entity_28481ebfc8
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      hw_tx => convert1_dout_net_x4,
      mac_io_phy_tx_phy_mode => phy_tx_phy_mode_net_x1,
      regtx_sw_tx_phy_mode => register26_q_net_x2,
      sw_tx => logical5_y_net_x2,
      phy_mode => mux_y_net_x0
    );

  pkt_buf_sel_412d479839: entity work.pkt_buf_sel_entity_412d479839
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      hw_tx => convert1_dout_net_x4,
      mac_io_phy_tx_pkt_buf => phy_tx_pkt_buf_net_x1,
      regtx_pkt_buf_sel => register15_q_net_x2,
      sw_tx => logical5_y_net_x2,
      pkt_buf => mux_y_net_x14
    );

  posedge1_95d3e0d45f: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      d => logical1_y_net_x1,
      q => logical1_y_net_x4
    );

  posedge2_6c78090f16: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      d => register2_q_net_x5,
      q => logical1_y_net_x6
    );

  posedge4_4c96bab1de: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      d => register1_q_net_x7,
      q => logical1_y_net_x2
    );

  posedge5_d5a0ca56ac: entity work.posedge1_entity_78541e5bea
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      d => logical1_y_net_x11,
      q => logical1_y_net_x3
    );

  register1: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x110,
      clk => clk_1_sg_x110,
      d => register4_q_net,
      en => "1",
      rst => "0",
      q => register1_q_net_x9
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x110,
      clk => clk_1_sg_x110,
      d(0) => register2_q_net_x0,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x8
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x110,
      clk => clk_1_sg_x110,
      d(0) => logical_y_net,
      en(0) => convert2_dout_net_x6,
      rst => "0",
      q(0) => register3_q_net_x9
    );

  register4: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x110,
      clk => clk_1_sg_x110,
      d => phy_tx_ant_mask_net_x0,
      en(0) => convert1_dout_net_x4,
      rst => "0",
      q => register4_q_net
    );

  rxen_control_677408d8f6: entity work.rxen_control_entity_677408d8f6
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      mac_tx_ant_mask => register1_q_net_x9,
      regtx_rc_rxen_enable => register1_q_net_x7,
      regtx_use_mac_ant_masks => register23_q_net_x5,
      rx => register2_q_net_x6,
      tx => register2_q_net_x9,
      rc_io_rxen => rc_rxen_x1,
      rc_io_txen_a => register5_q_net_x2,
      rc_io_txen_b => register1_q_net_x8,
      rc_io_txen_c => register2_q_net_x7,
      rc_io_txen_d => register3_q_net_x2
    );

  s_r_latch1_96bb620271: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      r => logical7_y_net_x0,
      s => logical4_y_net_x0,
      q => register2_q_net_x6
    );

  s_r_latch2_c31d9fc389: entity work.s_r_latch2_entity_c31d9fc389
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      r => logical8_y_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x0
    );

  s_r_latch_9c9835a519: entity work.s_r_latch1_entity_18268c34fe
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      r => logical6_y_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x9
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => mux_y_net_x0,
      y(0) => slice_y_net_x6
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => mux_y_net_x0,
      y(0) => slice1_y_net_x13
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => mux_y_net_x0,
      y(0) => slice2_y_net
    );

  tx_active_debug_signal_fb88e0bcc4: entity work.tx_active_debug_signal_entity_fb88e0bcc4
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      regtx_txrunning_output_sel => register24_q_net_x2,
      tx_active => register2_q_net_x5,
      register1_x0 => register1_q_net_x10
    );

  tx_gain_164a39bf58: entity work.tx_gain_entity_164a39bf58
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      hw_tx => convert1_dout_net_x4,
      phy_tx_gain_a => phy_tx_gain_a_net_x1,
      phy_tx_gain_b => phy_tx_gain_b_net_x1,
      phy_tx_gain_c => phy_tx_gain_c_net_x1,
      phy_tx_gain_d => phy_tx_gain_d_net_x1,
      sw_tx => logical5_y_net_x2,
      tx_gain_a => register1_q_net_x11,
      tx_gain_b => register3_q_net_x10,
      tx_gain_c => register5_q_net_x3,
      tx_gain_d => register7_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd"

entity wlan_phy_tx_pmd is
  port (
    axi_aresetn: in std_logic; 
    bram_din: in std_logic_vector(63 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_out: in std_logic_vector(31 downto 0); 
    data_out_x0: in std_logic_vector(31 downto 0); 
    data_out_x1: in std_logic_vector(31 downto 0); 
    data_out_x2: in std_logic_vector(31 downto 0); 
    data_out_x3: in std_logic_vector(31 downto 0); 
    data_out_x4: in std_logic_vector(31 downto 0); 
    data_out_x5: in std_logic_vector(31 downto 0); 
    dout: in std_logic_vector(31 downto 0); 
    dout_x0: in std_logic_vector(31 downto 0); 
    dout_x1: in std_logic_vector(31 downto 0); 
    dout_x2: in std_logic_vector(31 downto 0); 
    dout_x3: in std_logic_vector(31 downto 0); 
    dout_x4: in std_logic_vector(31 downto 0); 
    phy_tx_ant_mask: in std_logic_vector(3 downto 0); 
    phy_tx_gain_a: in std_logic_vector(5 downto 0); 
    phy_tx_gain_b: in std_logic_vector(5 downto 0); 
    phy_tx_gain_c: in std_logic_vector(5 downto 0); 
    phy_tx_gain_d: in std_logic_vector(5 downto 0); 
    phy_tx_phy_mode: in std_logic_vector(2 downto 0); 
    phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    phy_tx_start: in std_logic; 
    plb_ce_1: in std_logic; 
    plb_clk_1: in std_logic; 
    rc_phy_start: in std_logic; 
    s_axi_araddr: in std_logic_vector(31 downto 0); 
    s_axi_arburst: in std_logic_vector(1 downto 0); 
    s_axi_arcache: in std_logic_vector(3 downto 0); 
    s_axi_arid: in std_logic_vector(7 downto 0); 
    s_axi_arlen: in std_logic_vector(7 downto 0); 
    s_axi_arlock: in std_logic_vector(1 downto 0); 
    s_axi_arprot: in std_logic_vector(2 downto 0); 
    s_axi_arsize: in std_logic_vector(2 downto 0); 
    s_axi_arvalid: in std_logic; 
    s_axi_awaddr: in std_logic_vector(31 downto 0); 
    s_axi_awburst: in std_logic_vector(1 downto 0); 
    s_axi_awcache: in std_logic_vector(3 downto 0); 
    s_axi_awid: in std_logic_vector(7 downto 0); 
    s_axi_awlen: in std_logic_vector(7 downto 0); 
    s_axi_awlock: in std_logic_vector(1 downto 0); 
    s_axi_awprot: in std_logic_vector(2 downto 0); 
    s_axi_awsize: in std_logic_vector(2 downto 0); 
    s_axi_awvalid: in std_logic; 
    s_axi_bready: in std_logic; 
    s_axi_rready: in std_logic; 
    s_axi_wdata: in std_logic_vector(31 downto 0); 
    s_axi_wlast: in std_logic; 
    s_axi_wstrb: in std_logic_vector(3 downto 0); 
    s_axi_wvalid: in std_logic; 
    samp_ce: in std_logic; 
    bram_addr: out std_logic_vector(31 downto 0); 
    bram_dout: out std_logic_vector(63 downto 0); 
    bram_en: out std_logic; 
    bram_reset: out std_logic; 
    bram_wen: out std_logic_vector(7 downto 0); 
    data_in: out std_logic_vector(31 downto 0); 
    data_in_x0: out std_logic_vector(31 downto 0); 
    data_in_x1: out std_logic_vector(31 downto 0); 
    data_in_x2: out std_logic_vector(31 downto 0); 
    data_in_x3: out std_logic_vector(31 downto 0); 
    data_in_x4: out std_logic_vector(31 downto 0); 
    data_in_x5: out std_logic_vector(31 downto 0); 
    dbg_tx_running: out std_logic; 
    en: out std_logic; 
    en_x0: out std_logic; 
    en_x1: out std_logic; 
    en_x2: out std_logic; 
    en_x3: out std_logic; 
    en_x4: out std_logic; 
    en_x5: out std_logic; 
    phy_tx_done: out std_logic; 
    phy_tx_started: out std_logic; 
    rc_tx_gain_a: out std_logic_vector(5 downto 0); 
    rc_tx_gain_b: out std_logic_vector(5 downto 0); 
    rc_tx_gain_c: out std_logic_vector(5 downto 0); 
    rc_tx_gain_d: out std_logic_vector(5 downto 0); 
    rc_usr_rxen: out std_logic; 
    rc_usr_txen_a: out std_logic; 
    rc_usr_txen_b: out std_logic; 
    rc_usr_txen_c: out std_logic; 
    rc_usr_txen_d: out std_logic; 
    rfa_dac_i: out std_logic_vector(11 downto 0); 
    rfa_dac_q: out std_logic_vector(11 downto 0); 
    rfb_dac_i: out std_logic_vector(11 downto 0); 
    rfb_dac_q: out std_logic_vector(11 downto 0); 
    rfc_dac_i: out std_logic_vector(11 downto 0); 
    rfc_dac_q: out std_logic_vector(11 downto 0); 
    rfd_dac_i: out std_logic_vector(11 downto 0); 
    rfd_dac_q: out std_logic_vector(11 downto 0); 
    rx_sigs_invalid: out std_logic; 
    s_axi_arready: out std_logic; 
    s_axi_awready: out std_logic; 
    s_axi_bid: out std_logic_vector(7 downto 0); 
    s_axi_bresp: out std_logic_vector(1 downto 0); 
    s_axi_bvalid: out std_logic; 
    s_axi_rdata: out std_logic_vector(31 downto 0); 
    s_axi_rid: out std_logic_vector(7 downto 0); 
    s_axi_rlast: out std_logic; 
    s_axi_rresp: out std_logic_vector(1 downto 0); 
    s_axi_rvalid: out std_logic; 
    s_axi_wready: out std_logic
  );
end wlan_phy_tx_pmd;

architecture structural of wlan_phy_tx_pmd is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "wlan_phy_tx_pmd,sysgen_core,{black_box_isim_used=1,clock_period=6.25000000,clocking=Clock_Enables,sample_periods=1.00000000000 1.00000000000,testbench=0,total_blocks=2532,xilinx_accumulator_block=1,xilinx_adder_subtracter_block=13,xilinx_arithmetic_relational_operator_block=62,xilinx_assert_block=9,xilinx_axi_fifo_block_block=1,xilinx_bit_slice_extractor_block=203,xilinx_black_box_block=2,xilinx_bus_concatenator_block=35,xilinx_bus_multiplexer_block=57,xilinx_constant_block_block=156,xilinx_counter_block=16,xilinx_delay_block=72,xilinx_disregard_subsystem_for_generation_block=3,xilinx_dual_port_random_access_memory_block=2,xilinx_edk_core_block=1,xilinx_edk_processor_block=1,xilinx_fast_fourier_transform_8_0__block=1,xilinx_fifo_block_block=1,xilinx_gateway_in_block=37,xilinx_gateway_out_block=189,xilinx_inverter_block=56,xilinx_logical_block_block=170,xilinx_mcode_block_block=5,xilinx_multiplier_block=2,xilinx_register_block=138,xilinx_shared_memory_based_from_register_block=7,xilinx_shared_memory_based_to_register_block=7,xilinx_simulation_multiplexer_block=2,xilinx_single_port_read_only_memory_block=12,xilinx_system_generator_block=1,xilinx_type_converter_block=80,xilinx_type_reinterpreter_block=15,}";

  signal axi_aresetn_net: std_logic;
  signal axi_fifo_s_axis_tready_net_x5: std_logic;
  signal bram_addr_net: std_logic_vector(31 downto 0);
  signal bram_din_net: std_logic_vector(63 downto 0);
  signal bram_dout_net: std_logic_vector(63 downto 0);
  signal bram_en_net: std_logic;
  signal bram_reset_net: std_logic;
  signal bram_wen_net: std_logic_vector(7 downto 0);
  signal ce_1_sg_x111: std_logic;
  signal clk_1_sg_x111: std_logic;
  signal concat_y_net_x7: std_logic_vector(17 downto 0);
  signal convert1_dout_net_x4: std_logic;
  signal convert1_dout_net_x5: std_logic;
  signal convert2_dout_net_x1: std_logic;
  signal convert2_dout_net_x6: std_logic;
  signal data_in_net: std_logic_vector(31 downto 0);
  signal data_in_x0_net: std_logic_vector(31 downto 0);
  signal data_in_x1_net: std_logic_vector(31 downto 0);
  signal data_in_x2_net: std_logic_vector(31 downto 0);
  signal data_in_x3_net: std_logic_vector(31 downto 0);
  signal data_in_x4_net: std_logic_vector(31 downto 0);
  signal data_in_x5_net: std_logic_vector(31 downto 0);
  signal data_out_net: std_logic_vector(31 downto 0);
  signal data_out_x0_net: std_logic_vector(31 downto 0);
  signal data_out_x1_net: std_logic_vector(31 downto 0);
  signal data_out_x2_net: std_logic_vector(31 downto 0);
  signal data_out_x3_net: std_logic_vector(31 downto 0);
  signal data_out_x4_net: std_logic_vector(31 downto 0);
  signal data_out_x5_net: std_logic_vector(31 downto 0);
  signal dbg_tx_running_net: std_logic;
  signal delay1_q_net_x3: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay3_q_net_x3: std_logic;
  signal delay9_q_net_x3: std_logic;
  signal delay_q_net_x2: std_logic_vector(17 downto 0);
  signal delay_q_net_x8: std_logic;
  signal delay_q_net_x9: std_logic_vector(17 downto 0);
  signal dout_net: std_logic_vector(31 downto 0);
  signal dout_x0_net: std_logic_vector(31 downto 0);
  signal dout_x1_net: std_logic_vector(31 downto 0);
  signal dout_x2_net: std_logic_vector(31 downto 0);
  signal dout_x3_net: std_logic_vector(31 downto 0);
  signal dout_x4_net: std_logic_vector(31 downto 0);
  signal en_net: std_logic;
  signal en_x0_net: std_logic;
  signal en_x1_net: std_logic;
  signal en_x2_net: std_logic;
  signal en_x3_net: std_logic;
  signal en_x4_net: std_logic;
  signal en_x5_net: std_logic;
  signal fifo_dcount_net_x2: std_logic_vector(7 downto 0);
  signal i_x1: std_logic_vector(15 downto 0);
  signal iq_tlast_x1: std_logic;
  signal iq_tvalid_x1: std_logic;
  signal logical1_y_net_x13: std_logic;
  signal logical3_y_net_x7: std_logic;
  signal logical4_y_net_x7: std_logic;
  signal logical4_y_net_x9: std_logic;
  signal logical_y_net_x39: std_logic;
  signal mux1_y_net_x2: std_logic_vector(15 downto 0);
  signal mux2_y_net_x2: std_logic;
  signal mux3_y_net_x2: std_logic_vector(11 downto 0);
  signal mux3_y_net_x3: std_logic;
  signal mux4_y_net_x2: std_logic_vector(17 downto 0);
  signal mux4_y_net_x3: std_logic_vector(11 downto 0);
  signal mux6_y_net_x2: std_logic_vector(15 downto 0);
  signal mux_y_net_x14: std_logic_vector(3 downto 0);
  signal phy_tx_ant_mask_net: std_logic_vector(3 downto 0);
  signal phy_tx_done_net: std_logic;
  signal phy_tx_gain_a_net: std_logic_vector(5 downto 0);
  signal phy_tx_gain_b_net: std_logic_vector(5 downto 0);
  signal phy_tx_gain_c_net: std_logic_vector(5 downto 0);
  signal phy_tx_gain_d_net: std_logic_vector(5 downto 0);
  signal phy_tx_phy_mode_net: std_logic_vector(2 downto 0);
  signal phy_tx_pkt_buf_net: std_logic_vector(3 downto 0);
  signal phy_tx_start_net: std_logic;
  signal phy_tx_started_net: std_logic;
  signal plb_ce_1_sg_x1: std_logic;
  signal plb_clk_1_sg_x1: std_logic;
  signal q_x1: std_logic_vector(15 downto 0);
  signal rc_phy_start_net: std_logic;
  signal rc_tx_gain_a_net: std_logic_vector(5 downto 0);
  signal rc_tx_gain_b_net: std_logic_vector(5 downto 0);
  signal rc_tx_gain_c_net: std_logic_vector(5 downto 0);
  signal rc_tx_gain_d_net: std_logic_vector(5 downto 0);
  signal rc_usr_rxen_net: std_logic;
  signal rc_usr_txen_a_net: std_logic;
  signal rc_usr_txen_b_net: std_logic;
  signal rc_usr_txen_c_net: std_logic;
  signal rc_usr_txen_d_net: std_logic;
  signal register10_q_net_x2: std_logic_vector(5 downto 0);
  signal register11_q_net_x1: std_logic;
  signal register12_q_net_x1: std_logic;
  signal register13_q_net_x2: std_logic_vector(15 downto 0);
  signal register14_q_net_x2: std_logic_vector(15 downto 0);
  signal register15_q_net_x2: std_logic_vector(3 downto 0);
  signal register16_q_net_x3: std_logic_vector(7 downto 0);
  signal register17_q_net_x2: std_logic_vector(9 downto 0);
  signal register1_q_net_x7: std_logic;
  signal register1_q_net_x9: std_logic_vector(3 downto 0);
  signal register23_q_net_x5: std_logic;
  signal register24_q_net_x2: std_logic;
  signal register26_q_net_x2: std_logic_vector(2 downto 0);
  signal register27_q_net_x2: std_logic_vector(9 downto 0);
  signal register28_q_net_x2: std_logic_vector(9 downto 0);
  signal register2_q_net_x10: std_logic;
  signal register2_q_net_x6: std_logic;
  signal register3_q_net_x6: std_logic;
  signal register3_q_net_x9: std_logic;
  signal register4_q_net_x5: std_logic;
  signal register5_q_net_x5: std_logic;
  signal register6_q_net_x5: std_logic;
  signal register7_q_net_x2: std_logic;
  signal register8_q_net_x9: std_logic_vector(7 downto 0);
  signal register9_q_net_x3: std_logic_vector(7 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x6: std_logic_vector(15 downto 0);
  signal rfa_dac_i_net: std_logic_vector(11 downto 0);
  signal rfa_dac_q_net: std_logic_vector(11 downto 0);
  signal rfb_dac_i_net: std_logic_vector(11 downto 0);
  signal rfb_dac_q_net: std_logic_vector(11 downto 0);
  signal rfc_dac_i_net: std_logic_vector(11 downto 0);
  signal rfc_dac_q_net: std_logic_vector(11 downto 0);
  signal rfd_dac_i_net: std_logic_vector(11 downto 0);
  signal rfd_dac_q_net: std_logic_vector(11 downto 0);
  signal rx_sigs_invalid_net: std_logic;
  signal s_axi_araddr_net: std_logic_vector(31 downto 0);
  signal s_axi_arburst_net: std_logic_vector(1 downto 0);
  signal s_axi_arcache_net: std_logic_vector(3 downto 0);
  signal s_axi_arid_net: std_logic_vector(7 downto 0);
  signal s_axi_arlen_net: std_logic_vector(7 downto 0);
  signal s_axi_arlock_net: std_logic_vector(1 downto 0);
  signal s_axi_arprot_net: std_logic_vector(2 downto 0);
  signal s_axi_arready_net: std_logic;
  signal s_axi_arsize_net: std_logic_vector(2 downto 0);
  signal s_axi_arvalid_net: std_logic;
  signal s_axi_awaddr_net: std_logic_vector(31 downto 0);
  signal s_axi_awburst_net: std_logic_vector(1 downto 0);
  signal s_axi_awcache_net: std_logic_vector(3 downto 0);
  signal s_axi_awid_net: std_logic_vector(7 downto 0);
  signal s_axi_awlen_net: std_logic_vector(7 downto 0);
  signal s_axi_awlock_net: std_logic_vector(1 downto 0);
  signal s_axi_awprot_net: std_logic_vector(2 downto 0);
  signal s_axi_awready_net: std_logic;
  signal s_axi_awsize_net: std_logic_vector(2 downto 0);
  signal s_axi_awvalid_net: std_logic;
  signal s_axi_bid_net: std_logic_vector(7 downto 0);
  signal s_axi_bready_net: std_logic;
  signal s_axi_bresp_net: std_logic_vector(1 downto 0);
  signal s_axi_bvalid_net: std_logic;
  signal s_axi_rdata_net: std_logic_vector(31 downto 0);
  signal s_axi_rid_net: std_logic_vector(7 downto 0);
  signal s_axi_rlast_net: std_logic;
  signal s_axi_rready_net: std_logic;
  signal s_axi_rresp_net: std_logic_vector(1 downto 0);
  signal s_axi_rvalid_net: std_logic;
  signal s_axi_wdata_net: std_logic_vector(31 downto 0);
  signal s_axi_wlast_net: std_logic;
  signal s_axi_wready_net: std_logic;
  signal s_axi_wstrb_net: std_logic_vector(3 downto 0);
  signal s_axi_wvalid_net: std_logic;
  signal samp_ce_net: std_logic;
  signal slice1_y_net_x13: std_logic;
  signal slice_y_net_x6: std_logic;

begin
  axi_aresetn_net <= axi_aresetn;
  bram_din_net <= bram_din;
  ce_1_sg_x111 <= ce_1;
  clk_1_sg_x111 <= clk_1;
  data_out_net <= data_out;
  data_out_x0_net <= data_out_x0;
  data_out_x1_net <= data_out_x1;
  data_out_x2_net <= data_out_x2;
  data_out_x3_net <= data_out_x3;
  data_out_x4_net <= data_out_x4;
  data_out_x5_net <= data_out_x5;
  dout_net <= dout;
  dout_x0_net <= dout_x0;
  dout_x1_net <= dout_x1;
  dout_x2_net <= dout_x2;
  dout_x3_net <= dout_x3;
  dout_x4_net <= dout_x4;
  phy_tx_ant_mask_net <= phy_tx_ant_mask;
  phy_tx_gain_a_net <= phy_tx_gain_a;
  phy_tx_gain_b_net <= phy_tx_gain_b;
  phy_tx_gain_c_net <= phy_tx_gain_c;
  phy_tx_gain_d_net <= phy_tx_gain_d;
  phy_tx_phy_mode_net <= phy_tx_phy_mode;
  phy_tx_pkt_buf_net <= phy_tx_pkt_buf;
  phy_tx_start_net <= phy_tx_start;
  plb_ce_1_sg_x1 <= plb_ce_1;
  plb_clk_1_sg_x1 <= plb_clk_1;
  rc_phy_start_net <= rc_phy_start;
  s_axi_araddr_net <= s_axi_araddr;
  s_axi_arburst_net <= s_axi_arburst;
  s_axi_arcache_net <= s_axi_arcache;
  s_axi_arid_net <= s_axi_arid;
  s_axi_arlen_net <= s_axi_arlen;
  s_axi_arlock_net <= s_axi_arlock;
  s_axi_arprot_net <= s_axi_arprot;
  s_axi_arsize_net <= s_axi_arsize;
  s_axi_arvalid_net <= s_axi_arvalid;
  s_axi_awaddr_net <= s_axi_awaddr;
  s_axi_awburst_net <= s_axi_awburst;
  s_axi_awcache_net <= s_axi_awcache;
  s_axi_awid_net <= s_axi_awid;
  s_axi_awlen_net <= s_axi_awlen;
  s_axi_awlock_net <= s_axi_awlock;
  s_axi_awprot_net <= s_axi_awprot;
  s_axi_awsize_net <= s_axi_awsize;
  s_axi_awvalid_net <= s_axi_awvalid;
  s_axi_bready_net <= s_axi_bready;
  s_axi_rready_net <= s_axi_rready;
  s_axi_wdata_net <= s_axi_wdata;
  s_axi_wlast_net <= s_axi_wlast;
  s_axi_wstrb_net <= s_axi_wstrb;
  s_axi_wvalid_net <= s_axi_wvalid;
  samp_ce_net <= samp_ce;
  bram_addr <= bram_addr_net;
  bram_dout <= bram_dout_net;
  bram_en <= bram_en_net;
  bram_reset <= bram_reset_net;
  bram_wen <= bram_wen_net;
  data_in <= data_in_net;
  data_in_x0 <= data_in_x0_net;
  data_in_x1 <= data_in_x1_net;
  data_in_x2 <= data_in_x2_net;
  data_in_x3 <= data_in_x3_net;
  data_in_x4 <= data_in_x4_net;
  data_in_x5 <= data_in_x5_net;
  dbg_tx_running <= dbg_tx_running_net;
  en <= en_net;
  en_x0 <= en_x0_net;
  en_x1 <= en_x1_net;
  en_x2 <= en_x2_net;
  en_x3 <= en_x3_net;
  en_x4 <= en_x4_net;
  en_x5 <= en_x5_net;
  phy_tx_done <= phy_tx_done_net;
  phy_tx_started <= phy_tx_started_net;
  rc_tx_gain_a <= rc_tx_gain_a_net;
  rc_tx_gain_b <= rc_tx_gain_b_net;
  rc_tx_gain_c <= rc_tx_gain_c_net;
  rc_tx_gain_d <= rc_tx_gain_d_net;
  rc_usr_rxen <= rc_usr_rxen_net;
  rc_usr_txen_a <= rc_usr_txen_a_net;
  rc_usr_txen_b <= rc_usr_txen_b_net;
  rc_usr_txen_c <= rc_usr_txen_c_net;
  rc_usr_txen_d <= rc_usr_txen_d_net;
  rfa_dac_i <= rfa_dac_i_net;
  rfa_dac_q <= rfa_dac_q_net;
  rfb_dac_i <= rfb_dac_i_net;
  rfb_dac_q <= rfb_dac_q_net;
  rfc_dac_i <= rfc_dac_i_net;
  rfc_dac_q <= rfc_dac_q_net;
  rfd_dac_i <= rfd_dac_i_net;
  rfd_dac_q <= rfd_dac_q_net;
  rx_sigs_invalid <= rx_sigs_invalid_net;
  s_axi_arready <= s_axi_arready_net;
  s_axi_awready <= s_axi_awready_net;
  s_axi_bid <= s_axi_bid_net;
  s_axi_bresp <= s_axi_bresp_net;
  s_axi_bvalid <= s_axi_bvalid_net;
  s_axi_rdata <= s_axi_rdata_net;
  s_axi_rid <= s_axi_rid_net;
  s_axi_rlast <= s_axi_rlast_net;
  s_axi_rresp <= s_axi_rresp_net;
  s_axi_rvalid <= s_axi_rvalid_net;
  s_axi_wready <= s_axi_wready_net;

  edk_processor_de00edcbbe: entity work.edk_processor_entity_de00edcbbe
    port map (
      axi_aresetn => axi_aresetn_net,
      from_register => data_out_net,
      plb_ce_1 => plb_ce_1_sg_x1,
      plb_clk_1 => plb_clk_1_sg_x1,
      s_axi_araddr => s_axi_araddr_net,
      s_axi_arburst => s_axi_arburst_net,
      s_axi_arcache => s_axi_arcache_net,
      s_axi_arid => s_axi_arid_net,
      s_axi_arlen => s_axi_arlen_net,
      s_axi_arlock => s_axi_arlock_net,
      s_axi_arprot => s_axi_arprot_net,
      s_axi_arsize => s_axi_arsize_net,
      s_axi_arvalid => s_axi_arvalid_net,
      s_axi_awaddr => s_axi_awaddr_net,
      s_axi_awburst => s_axi_awburst_net,
      s_axi_awcache => s_axi_awcache_net,
      s_axi_awid => s_axi_awid_net,
      s_axi_awlen => s_axi_awlen_net,
      s_axi_awlock => s_axi_awlock_net,
      s_axi_awprot => s_axi_awprot_net,
      s_axi_awsize => s_axi_awsize_net,
      s_axi_awvalid => s_axi_awvalid_net,
      s_axi_bready => s_axi_bready_net,
      s_axi_rready => s_axi_rready_net,
      s_axi_wdata => s_axi_wdata_net,
      s_axi_wlast => s_axi_wlast_net,
      s_axi_wstrb => s_axi_wstrb_net,
      s_axi_wvalid => s_axi_wvalid_net,
      to_register => dout_net,
      to_register1 => dout_x0_net,
      to_register2 => dout_x1_net,
      to_register3 => dout_x2_net,
      to_register4 => dout_x3_net,
      to_register5 => dout_x4_net,
      memmap_x0 => s_axi_arready_net,
      memmap_x1 => s_axi_awready_net,
      memmap_x10 => s_axi_wready_net,
      memmap_x11 => data_in_net,
      memmap_x12 => en_net,
      memmap_x13 => data_in_x0_net,
      memmap_x14 => en_x0_net,
      memmap_x15 => data_in_x1_net,
      memmap_x16 => en_x1_net,
      memmap_x17 => data_in_x2_net,
      memmap_x18 => en_x2_net,
      memmap_x19 => data_in_x3_net,
      memmap_x2 => s_axi_bid_net,
      memmap_x20 => en_x3_net,
      memmap_x21 => data_in_x4_net,
      memmap_x22 => en_x4_net,
      memmap_x3 => s_axi_bresp_net,
      memmap_x4 => s_axi_bvalid_net,
      memmap_x5 => s_axi_rdata_net,
      memmap_x6 => s_axi_rid_net,
      memmap_x7 => s_axi_rlast_net,
      memmap_x8 => s_axi_rresp_net,
      memmap_x9 => s_axi_rvalid_net
    );

  ht_preamble_gen_624eef30fb: entity work.ht_preamble_gen_entity_624eef30fb
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      iq_fifo_tready => axi_fifo_s_axis_tready_net_x5,
      start => logical4_y_net_x7,
      sym_cfg => concat_y_net_x7,
      tx_reset => logical_y_net_x39,
      delay1_x0 => iq_tvalid_x1,
      delay2_x0 => iq_tlast_x1,
      ht_training_q_x0 => q_x1,
      iq_stream => i_x1,
      sym_cfg_x0 => delay_q_net_x2
    );

  ifft_and_cyclic_prefix_d9041c6806: entity work.ifft_and_cyclic_prefix_entity_d9041c6806
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      i => mux6_y_net_x2,
      iq_tlast => mux3_y_net_x3,
      iq_valid => mux2_y_net_x2,
      logical => logical_y_net_x39,
      q => mux1_y_net_x2,
      register10 => register10_q_net_x2,
      register8 => register8_q_net_x9,
      register9 => register9_q_net_x3,
      sym_cfg => mux4_y_net_x2,
      fifo_tready => axi_fifo_s_axis_tready_net_x5,
      i_x0 => reinterpret2_output_port_net_x6,
      iq_valid_x0 => delay3_q_net_x3,
      q_x0 => reinterpret3_output_port_net_x6
    );

  mux_e0e38b1125: entity work.mux_entity_e0e38b1125
    port map (
      delay => delay_q_net_x8,
      delay1 => delay1_q_net_x3,
      ht_preamble_gen => iq_tvalid_x1,
      ht_preamble_gen_x0 => iq_tlast_x1,
      ht_preamble_gen_x1 => q_x1,
      mux4_x0 => mux4_y_net_x3,
      preamble_iq => i_x1,
      preamble_sym_cfg => delay_q_net_x2,
      psdu_iq => mux3_y_net_x2,
      psdu_sym_cfg => delay_q_net_x9,
      i => mux6_y_net_x2,
      iq_tlast => mux3_y_net_x3,
      iq_tvalid => mux2_y_net_x2,
      q => mux1_y_net_x2,
      sym_cfg => mux4_y_net_x2
    );

  ofdm_symbol_ctrl_c16241a486: entity work.ofdm_symbol_ctrl_entity_c16241a486
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      convert2 => convert2_dout_net_x6,
      data_done => delay9_q_net_x3,
      logical3_x0 => logical3_y_net_x7,
      output_fifo_occ => fifo_dcount_net_x2,
      register8 => register8_q_net_x9,
      slice => slice_y_net_x6,
      slice1 => slice1_y_net_x13,
      start_tx => register3_q_net_x9,
      sym_done => mux3_y_net_x3,
      tx_reset => logical_y_net_x39,
      start_sym => logical4_y_net_x7,
      sym_cfg => concat_y_net_x7
    );

  preamble_outputs_82fcc722dc: entity work.\preamble___outputs_entity_82fcc722dc\
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      i => reinterpret2_output_port_net_x6,
      iq_tvalid => delay3_q_net_x3,
      q => reinterpret3_output_port_net_x6,
      register1 => register1_q_net_x9,
      register13 => register13_q_net_x2,
      register14 => register14_q_net_x2,
      register23 => register23_q_net_x5,
      register3_x0 => register3_q_net_x6,
      register4_x0 => register4_q_net_x5,
      register5 => register5_q_net_x5,
      register6 => register6_q_net_x5,
      tx_iq_samp_ce => convert2_dout_net_x6,
      tx_reset => logical_y_net_x39,
      tx_start => register3_q_net_x9,
      dac_outputs => rfa_dac_i_net,
      dac_outputs_x0 => rfa_dac_q_net,
      dac_outputs_x1 => rfb_dac_i_net,
      dac_outputs_x2 => rfb_dac_q_net,
      dac_outputs_x3 => rfc_dac_i_net,
      dac_outputs_x4 => rfc_dac_q_net,
      dac_outputs_x5 => rfd_dac_i_net,
      dac_outputs_x6 => rfd_dac_q_net,
      fifo => fifo_dcount_net_x2,
      last_samp_output_to_dacs => delay2_q_net_x1
    );

  psdu_syms_gen_1449f55c9b: entity work.psdu_syms_gen_entity_1449f55c9b
    port map (
      bram_din => bram_din_net,
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      iq_fifo_tready => axi_fifo_s_axis_tready_net_x5,
      logical => logical_y_net_x39,
      logical3 => logical3_y_net_x7,
      mux => mux_y_net_x14,
      register16 => register16_q_net_x3,
      register2 => register2_q_net_x6,
      register8 => register8_q_net_x9,
      slice => slice_y_net_x6,
      slice1 => slice1_y_net_x13,
      start_sym => logical4_y_net_x7,
      sym_cfg => concat_y_net_x7,
      data_done => delay9_q_net_x3,
      iq_stream => mux3_y_net_x2,
      modulate => delay_q_net_x8,
      modulate_x0 => delay1_q_net_x3,
      modulate_x1 => mux4_y_net_x3,
      pkt_data => bram_addr_net,
      pkt_data_x0 => bram_en_net,
      pkt_data_x1 => bram_reset_net,
      pkt_data_x2 => bram_dout_net,
      pkt_data_x3 => bram_wen_net,
      pkt_data_x4 => logical4_y_net_x9,
      sym_cfg_x0 => delay_q_net_x9
    );

  radio_controller_mac_io_c70eccdf43: entity work.\radio_controller___mac_io_entity_c70eccdf43\
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      phy_tx_start => phy_tx_start_net,
      rc_phy_start => rc_phy_start_net,
      mac_io_phy_tx_start => convert1_dout_net_x4,
      rc_io_phy_start => convert2_dout_net_x1
    );

  registers_2d8965b1e5: entity work.registers_entity_2d8965b1e5
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      from_register1 => data_out_x0_net,
      from_register2 => data_out_x1_net,
      from_register3 => data_out_x2_net,
      from_register4 => data_out_x3_net,
      from_register5 => data_out_x4_net,
      from_register6 => data_out_x5_net,
      register2_x0 => register2_q_net_x10,
      constant_x1 => en_x5_net,
      register20_x0 => data_in_x5_net,
      regtx_anta_tx_en => register3_q_net_x6,
      regtx_antb_tx_en => register4_q_net_x5,
      regtx_antc_tx_en => register5_q_net_x5,
      regtx_antd_tx_en => register6_q_net_x5,
      regtx_cp_len => register9_q_net_x3,
      regtx_fft_scaling => register10_q_net_x2,
      regtx_num_sc => register8_q_net_x9,
      regtx_pkt_buf_addr_offset => register16_q_net_x3,
      regtx_pkt_buf_sel => register15_q_net_x2,
      regtx_posttx_extension => register17_q_net_x2,
      regtx_posttx_rf_en_extension => register27_q_net_x2,
      regtx_posttx_rxsig_valid => register28_q_net_x2,
      regtx_rc_rxen_enable => register1_q_net_x7,
      regtx_reset => register7_q_net_x2,
      regtx_reset_scrambling_lfsr_perpkt => register2_q_net_x6,
      regtx_scaling_payload => register14_q_net_x2,
      regtx_scaling_preamble => register13_q_net_x2,
      regtx_start_direct => register11_q_net_x1,
      regtx_start_indirect => register12_q_net_x1,
      regtx_sw_tx_phy_mode => register26_q_net_x2,
      regtx_txrunning_output_sel => register24_q_net_x2,
      regtx_use_mac_ant_masks => register23_q_net_x5
    );

  resets_24d0a1b807: entity work.resets_entity_24d0a1b807
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      last_samp_output_to_dacs => delay2_q_net_x1,
      regtx_reset => register7_q_net_x2,
      tx_sig_decode_error => logical4_y_net_x9,
      tx_force_reset => convert1_dout_net_x5,
      tx_phy_done => logical1_y_net_x13,
      tx_reset => logical_y_net_x39
    );

  sampling_clock_a1a467035e: entity work.sampling_clock_entity_a1a467035e
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      samp_ce => samp_ce_net,
      tx_iq_samp_ce => convert2_dout_net_x6
    );

  start_ctrl_3ba2a032ad: entity work.start_ctrl_entity_3ba2a032ad
    port map (
      ce_1 => ce_1_sg_x111,
      clk_1 => clk_1_sg_x111,
      mac_io_phy_tx_ant_mask => phy_tx_ant_mask_net,
      mac_io_phy_tx_start => convert1_dout_net_x4,
      phy_tx_gain_a => phy_tx_gain_a_net,
      phy_tx_gain_b => phy_tx_gain_b_net,
      phy_tx_gain_c => phy_tx_gain_c_net,
      phy_tx_gain_d => phy_tx_gain_d_net,
      phy_tx_phy_mode => phy_tx_phy_mode_net,
      phy_tx_pkt_buf => phy_tx_pkt_buf_net,
      rc_io_phy_start => convert2_dout_net_x1,
      registers => register15_q_net_x2,
      registers_x0 => register17_q_net_x2,
      registers_x1 => register23_q_net_x5,
      registers_x2 => register24_q_net_x2,
      registers_x3 => register26_q_net_x2,
      registers_x4 => register27_q_net_x2,
      registers_x5 => register28_q_net_x2,
      regtx_rc_rxen_enable => register1_q_net_x7,
      regtx_start_direct => register11_q_net_x1,
      regtx_start_indirect => register12_q_net_x1,
      tx_force_reset => convert1_dout_net_x5,
      tx_iq_samp_ce => convert2_dout_net_x6,
      tx_phy_done => logical1_y_net_x13,
      mac_io_phy_tx_done => phy_tx_done_net,
      mac_io_phy_tx_started => phy_tx_started_net,
      mac_tx_ant_mask => register1_q_net_x9,
      phy_start => register3_q_net_x9,
      rc_io_tx_gain_a => rc_tx_gain_a_net,
      rc_io_tx_gain_b => rc_tx_gain_b_net,
      rc_io_tx_gain_c => rc_tx_gain_c_net,
      rc_io_tx_gain_d => rc_tx_gain_d_net,
      register2_x0 => rx_sigs_invalid_net,
      regtx_tx_running => register2_q_net_x10,
      rxen_control => rc_usr_txen_b_net,
      rxen_control_x0 => rc_usr_txen_c_net,
      rxen_control_x1 => rc_usr_txen_d_net,
      rxen_control_x2 => rc_usr_rxen_net,
      rxen_control_x3 => rc_usr_txen_a_net,
      tx_active_debug_signal => dbg_tx_running_net,
      tx_phy_mode_11ag => slice_y_net_x6,
      tx_phy_mode_11n => slice1_y_net_x13,
      tx_phy_mode_11n_ac => logical3_y_net_x7,
      tx_pkt_buf_sel => mux_y_net_x14
    );

end structural;
